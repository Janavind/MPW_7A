VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 420.740 800.600 421.060 800.660 ;
        RECT 2901.290 800.600 2901.610 800.660 ;
        RECT 420.740 800.460 2901.610 800.600 ;
        RECT 420.740 800.400 421.060 800.460 ;
        RECT 2901.290 800.400 2901.610 800.460 ;
      LAYER via ;
        RECT 420.770 800.400 421.030 800.660 ;
        RECT 2901.320 800.400 2901.580 800.660 ;
      LAYER met2 ;
        RECT 420.770 800.370 421.030 800.690 ;
        RECT 2901.320 800.370 2901.580 800.690 ;
        RECT 420.830 800.000 420.970 800.370 ;
        RECT 420.790 796.000 421.070 800.000 ;
        RECT 2901.380 33.165 2901.520 800.370 ;
        RECT 2901.310 32.795 2901.590 33.165 ;
      LAYER via2 ;
        RECT 2901.310 32.840 2901.590 33.120 ;
      LAYER met3 ;
        RECT 2901.285 33.130 2901.615 33.145 ;
        RECT 2917.600 33.130 2924.800 33.580 ;
        RECT 2901.285 32.830 2924.800 33.130 ;
        RECT 2901.285 32.815 2901.615 32.830 ;
        RECT 2917.600 32.380 2924.800 32.830 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 489.970 2284.020 490.290 2284.080 ;
        RECT 2900.830 2284.020 2901.150 2284.080 ;
        RECT 489.970 2283.880 2901.150 2284.020 ;
        RECT 489.970 2283.820 490.290 2283.880 ;
        RECT 2900.830 2283.820 2901.150 2283.880 ;
      LAYER via ;
        RECT 490.000 2283.820 490.260 2284.080 ;
        RECT 2900.860 2283.820 2901.120 2284.080 ;
      LAYER met2 ;
        RECT 2900.850 2290.395 2901.130 2290.765 ;
        RECT 2900.920 2284.110 2901.060 2290.395 ;
        RECT 490.000 2283.790 490.260 2284.110 ;
        RECT 2900.860 2283.790 2901.120 2284.110 ;
        RECT 490.060 800.000 490.200 2283.790 ;
        RECT 489.790 799.270 490.200 800.000 ;
        RECT 489.790 796.000 490.070 799.270 ;
      LAYER via2 ;
        RECT 2900.850 2290.440 2901.130 2290.720 ;
      LAYER met3 ;
        RECT 2900.825 2290.730 2901.155 2290.745 ;
        RECT 2917.600 2290.730 2924.800 2291.180 ;
        RECT 2900.825 2290.430 2924.800 2290.730 ;
        RECT 2900.825 2290.415 2901.155 2290.430 ;
        RECT 2917.600 2289.980 2924.800 2290.430 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.870 2553.300 497.190 2553.360 ;
        RECT 2900.830 2553.300 2901.150 2553.360 ;
        RECT 496.870 2553.160 2901.150 2553.300 ;
        RECT 496.870 2553.100 497.190 2553.160 ;
        RECT 2900.830 2553.100 2901.150 2553.160 ;
      LAYER via ;
        RECT 496.900 2553.100 497.160 2553.360 ;
        RECT 2900.860 2553.100 2901.120 2553.360 ;
      LAYER met2 ;
        RECT 2900.850 2556.275 2901.130 2556.645 ;
        RECT 2900.920 2553.390 2901.060 2556.275 ;
        RECT 496.900 2553.070 497.160 2553.390 ;
        RECT 2900.860 2553.070 2901.120 2553.390 ;
        RECT 496.960 800.000 497.100 2553.070 ;
        RECT 496.690 799.270 497.100 800.000 ;
        RECT 496.690 796.000 496.970 799.270 ;
      LAYER via2 ;
        RECT 2900.850 2556.320 2901.130 2556.600 ;
      LAYER met3 ;
        RECT 2900.825 2556.610 2901.155 2556.625 ;
        RECT 2917.600 2556.610 2924.800 2557.060 ;
        RECT 2900.825 2556.310 2924.800 2556.610 ;
        RECT 2900.825 2556.295 2901.155 2556.310 ;
        RECT 2917.600 2555.860 2924.800 2556.310 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 503.770 2815.440 504.090 2815.500 ;
        RECT 2898.990 2815.440 2899.310 2815.500 ;
        RECT 503.770 2815.300 2899.310 2815.440 ;
        RECT 503.770 2815.240 504.090 2815.300 ;
        RECT 2898.990 2815.240 2899.310 2815.300 ;
      LAYER via ;
        RECT 503.800 2815.240 504.060 2815.500 ;
        RECT 2899.020 2815.240 2899.280 2815.500 ;
      LAYER met2 ;
        RECT 2899.010 2821.475 2899.290 2821.845 ;
        RECT 2899.080 2815.530 2899.220 2821.475 ;
        RECT 503.800 2815.210 504.060 2815.530 ;
        RECT 2899.020 2815.210 2899.280 2815.530 ;
        RECT 503.860 800.000 504.000 2815.210 ;
        RECT 503.590 799.270 504.000 800.000 ;
        RECT 503.590 796.000 503.870 799.270 ;
      LAYER via2 ;
        RECT 2899.010 2821.520 2899.290 2821.800 ;
      LAYER met3 ;
        RECT 2898.985 2821.810 2899.315 2821.825 ;
        RECT 2917.600 2821.810 2924.800 2822.260 ;
        RECT 2898.985 2821.510 2924.800 2821.810 ;
        RECT 2898.985 2821.495 2899.315 2821.510 ;
        RECT 2917.600 2821.060 2924.800 2821.510 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.670 3084.380 510.990 3084.440 ;
        RECT 2900.830 3084.380 2901.150 3084.440 ;
        RECT 510.670 3084.240 2901.150 3084.380 ;
        RECT 510.670 3084.180 510.990 3084.240 ;
        RECT 2900.830 3084.180 2901.150 3084.240 ;
      LAYER via ;
        RECT 510.700 3084.180 510.960 3084.440 ;
        RECT 2900.860 3084.180 2901.120 3084.440 ;
      LAYER met2 ;
        RECT 2900.850 3087.355 2901.130 3087.725 ;
        RECT 2900.920 3084.470 2901.060 3087.355 ;
        RECT 510.700 3084.150 510.960 3084.470 ;
        RECT 2900.860 3084.150 2901.120 3084.470 ;
        RECT 510.760 800.000 510.900 3084.150 ;
        RECT 510.490 799.270 510.900 800.000 ;
        RECT 510.490 796.000 510.770 799.270 ;
      LAYER via2 ;
        RECT 2900.850 3087.400 2901.130 3087.680 ;
      LAYER met3 ;
        RECT 2900.825 3087.690 2901.155 3087.705 ;
        RECT 2917.600 3087.690 2924.800 3088.140 ;
        RECT 2900.825 3087.390 2924.800 3087.690 ;
        RECT 2900.825 3087.375 2901.155 3087.390 ;
        RECT 2917.600 3086.940 2924.800 3087.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.570 3353.660 517.890 3353.720 ;
        RECT 2900.830 3353.660 2901.150 3353.720 ;
        RECT 517.570 3353.520 2901.150 3353.660 ;
        RECT 517.570 3353.460 517.890 3353.520 ;
        RECT 2900.830 3353.460 2901.150 3353.520 ;
      LAYER via ;
        RECT 517.600 3353.460 517.860 3353.720 ;
        RECT 2900.860 3353.460 2901.120 3353.720 ;
      LAYER met2 ;
        RECT 517.600 3353.430 517.860 3353.750 ;
        RECT 2900.860 3353.605 2901.120 3353.750 ;
        RECT 517.660 800.000 517.800 3353.430 ;
        RECT 2900.850 3353.235 2901.130 3353.605 ;
        RECT 517.390 799.270 517.800 800.000 ;
        RECT 517.390 796.000 517.670 799.270 ;
      LAYER via2 ;
        RECT 2900.850 3353.280 2901.130 3353.560 ;
      LAYER met3 ;
        RECT 2900.825 3353.570 2901.155 3353.585 ;
        RECT 2917.600 3353.570 2924.800 3354.020 ;
        RECT 2900.825 3353.270 2924.800 3353.570 ;
        RECT 2900.825 3353.255 2901.155 3353.270 ;
        RECT 2917.600 3352.820 2924.800 3353.270 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.470 817.600 524.790 817.660 ;
        RECT 2794.570 817.600 2794.890 817.660 ;
        RECT 524.470 817.460 2794.890 817.600 ;
        RECT 524.470 817.400 524.790 817.460 ;
        RECT 2794.570 817.400 2794.890 817.460 ;
      LAYER via ;
        RECT 524.500 817.400 524.760 817.660 ;
        RECT 2794.600 817.400 2794.860 817.660 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3512.170 2798.480 3517.600 ;
        RECT 2794.660 3512.030 2798.480 3512.170 ;
        RECT 2794.660 817.690 2794.800 3512.030 ;
        RECT 524.500 817.370 524.760 817.690 ;
        RECT 2794.600 817.370 2794.860 817.690 ;
        RECT 524.560 800.000 524.700 817.370 ;
        RECT 524.290 799.270 524.700 800.000 ;
        RECT 524.290 796.000 524.570 799.270 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.370 817.940 531.690 818.000 ;
        RECT 2470.270 817.940 2470.590 818.000 ;
        RECT 531.370 817.800 2470.590 817.940 ;
        RECT 531.370 817.740 531.690 817.800 ;
        RECT 2470.270 817.740 2470.590 817.800 ;
      LAYER via ;
        RECT 531.400 817.740 531.660 818.000 ;
        RECT 2470.300 817.740 2470.560 818.000 ;
      LAYER met2 ;
        RECT 2470.360 3517.910 2473.260 3518.050 ;
        RECT 2470.360 818.030 2470.500 3517.910 ;
        RECT 2473.120 3517.370 2473.260 3517.910 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2473.120 3517.230 2474.180 3517.370 ;
        RECT 531.400 817.710 531.660 818.030 ;
        RECT 2470.300 817.710 2470.560 818.030 ;
        RECT 531.460 800.000 531.600 817.710 ;
        RECT 531.190 799.270 531.600 800.000 ;
        RECT 531.190 796.000 531.470 799.270 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.270 818.280 538.590 818.340 ;
        RECT 2145.970 818.280 2146.290 818.340 ;
        RECT 538.270 818.140 2146.290 818.280 ;
        RECT 538.270 818.080 538.590 818.140 ;
        RECT 2145.970 818.080 2146.290 818.140 ;
      LAYER via ;
        RECT 538.300 818.080 538.560 818.340 ;
        RECT 2146.000 818.080 2146.260 818.340 ;
      LAYER met2 ;
        RECT 2146.060 3517.910 2148.500 3518.050 ;
        RECT 2146.060 818.370 2146.200 3517.910 ;
        RECT 2148.360 3517.370 2148.500 3517.910 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3517.370 2149.420 3517.600 ;
        RECT 2148.360 3517.230 2149.420 3517.370 ;
        RECT 538.300 818.050 538.560 818.370 ;
        RECT 2146.000 818.050 2146.260 818.370 ;
        RECT 538.360 800.000 538.500 818.050 ;
        RECT 538.090 799.270 538.500 800.000 ;
        RECT 538.090 796.000 538.370 799.270 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.170 818.620 545.490 818.680 ;
        RECT 1821.670 818.620 1821.990 818.680 ;
        RECT 545.170 818.480 1821.990 818.620 ;
        RECT 545.170 818.420 545.490 818.480 ;
        RECT 1821.670 818.420 1821.990 818.480 ;
      LAYER via ;
        RECT 545.200 818.420 545.460 818.680 ;
        RECT 1821.700 818.420 1821.960 818.680 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3512.170 1825.120 3517.600 ;
        RECT 1821.760 3512.030 1825.120 3512.170 ;
        RECT 1821.760 818.710 1821.900 3512.030 ;
        RECT 545.200 818.390 545.460 818.710 ;
        RECT 1821.700 818.390 1821.960 818.710 ;
        RECT 545.260 800.000 545.400 818.390 ;
        RECT 544.990 799.270 545.400 800.000 ;
        RECT 544.990 796.000 545.270 799.270 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.070 818.960 552.390 819.020 ;
        RECT 1497.370 818.960 1497.690 819.020 ;
        RECT 552.070 818.820 1497.690 818.960 ;
        RECT 552.070 818.760 552.390 818.820 ;
        RECT 1497.370 818.760 1497.690 818.820 ;
      LAYER via ;
        RECT 552.100 818.760 552.360 819.020 ;
        RECT 1497.400 818.760 1497.660 819.020 ;
      LAYER met2 ;
        RECT 1497.460 3517.910 1499.900 3518.050 ;
        RECT 1497.460 819.050 1497.600 3517.910 ;
        RECT 1499.760 3517.370 1499.900 3517.910 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3517.370 1500.820 3517.600 ;
        RECT 1499.760 3517.230 1500.820 3517.370 ;
        RECT 552.100 818.730 552.360 819.050 ;
        RECT 1497.400 818.730 1497.660 819.050 ;
        RECT 552.160 800.000 552.300 818.730 ;
        RECT 551.890 799.270 552.300 800.000 ;
        RECT 551.890 796.000 552.170 799.270 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 429.250 800.940 429.570 801.000 ;
        RECT 2902.210 800.940 2902.530 801.000 ;
        RECT 429.250 800.800 2902.530 800.940 ;
        RECT 429.250 800.740 429.570 800.800 ;
        RECT 2902.210 800.740 2902.530 800.800 ;
      LAYER via ;
        RECT 429.280 800.740 429.540 801.000 ;
        RECT 2902.240 800.740 2902.500 801.000 ;
      LAYER met2 ;
        RECT 429.280 800.710 429.540 801.030 ;
        RECT 2902.240 800.710 2902.500 801.030 ;
        RECT 427.690 799.410 427.970 800.000 ;
        RECT 429.340 799.410 429.480 800.710 ;
        RECT 427.690 799.270 429.480 799.410 ;
        RECT 427.690 796.000 427.970 799.270 ;
        RECT 2902.300 231.725 2902.440 800.710 ;
        RECT 2902.230 231.355 2902.510 231.725 ;
      LAYER via2 ;
        RECT 2902.230 231.400 2902.510 231.680 ;
      LAYER met3 ;
        RECT 2902.205 231.690 2902.535 231.705 ;
        RECT 2917.600 231.690 2924.800 232.140 ;
        RECT 2902.205 231.390 2924.800 231.690 ;
        RECT 2902.205 231.375 2902.535 231.390 ;
        RECT 2917.600 230.940 2924.800 231.390 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.970 819.300 559.290 819.360 ;
        RECT 1173.070 819.300 1173.390 819.360 ;
        RECT 558.970 819.160 1173.390 819.300 ;
        RECT 558.970 819.100 559.290 819.160 ;
        RECT 1173.070 819.100 1173.390 819.160 ;
      LAYER via ;
        RECT 559.000 819.100 559.260 819.360 ;
        RECT 1173.100 819.100 1173.360 819.360 ;
      LAYER met2 ;
        RECT 1173.160 3517.910 1175.140 3518.050 ;
        RECT 1173.160 819.390 1173.300 3517.910 ;
        RECT 1175.000 3517.370 1175.140 3517.910 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3517.370 1176.060 3517.600 ;
        RECT 1175.000 3517.230 1176.060 3517.370 ;
        RECT 559.000 819.070 559.260 819.390 ;
        RECT 1173.100 819.070 1173.360 819.390 ;
        RECT 559.060 800.000 559.200 819.070 ;
        RECT 558.790 799.270 559.200 800.000 ;
        RECT 558.790 796.000 559.070 799.270 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 565.870 826.440 566.190 826.500 ;
        RECT 848.770 826.440 849.090 826.500 ;
        RECT 565.870 826.300 849.090 826.440 ;
        RECT 565.870 826.240 566.190 826.300 ;
        RECT 848.770 826.240 849.090 826.300 ;
      LAYER via ;
        RECT 565.900 826.240 566.160 826.500 ;
        RECT 848.800 826.240 849.060 826.500 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3512.170 851.760 3517.600 ;
        RECT 848.860 3512.030 851.760 3512.170 ;
        RECT 848.860 826.530 849.000 3512.030 ;
        RECT 565.900 826.210 566.160 826.530 ;
        RECT 848.800 826.210 849.060 826.530 ;
        RECT 565.960 800.000 566.100 826.210 ;
        RECT 565.690 799.270 566.100 800.000 ;
        RECT 565.690 796.000 565.970 799.270 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.470 819.640 524.790 819.700 ;
        RECT 572.770 819.640 573.090 819.700 ;
        RECT 524.470 819.500 573.090 819.640 ;
        RECT 524.470 819.440 524.790 819.500 ;
        RECT 572.770 819.440 573.090 819.500 ;
      LAYER via ;
        RECT 524.500 819.440 524.760 819.700 ;
        RECT 572.800 819.440 573.060 819.700 ;
      LAYER met2 ;
        RECT 524.560 3517.910 526.540 3518.050 ;
        RECT 524.560 819.730 524.700 3517.910 ;
        RECT 526.400 3517.370 526.540 3517.910 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3517.370 527.460 3517.600 ;
        RECT 526.400 3517.230 527.460 3517.370 ;
        RECT 524.500 819.410 524.760 819.730 ;
        RECT 572.800 819.410 573.060 819.730 ;
        RECT 572.860 800.000 573.000 819.410 ;
        RECT 572.590 799.270 573.000 800.000 ;
        RECT 572.590 796.000 572.870 799.270 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 200.170 826.100 200.490 826.160 ;
        RECT 579.670 826.100 579.990 826.160 ;
        RECT 200.170 825.960 579.990 826.100 ;
        RECT 200.170 825.900 200.490 825.960 ;
        RECT 579.670 825.900 579.990 825.960 ;
      LAYER via ;
        RECT 200.200 825.900 200.460 826.160 ;
        RECT 579.700 825.900 579.960 826.160 ;
      LAYER met2 ;
        RECT 200.260 3517.910 201.780 3518.050 ;
        RECT 200.260 826.190 200.400 3517.910 ;
        RECT 201.640 3517.370 201.780 3517.910 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3517.370 202.700 3517.600 ;
        RECT 201.640 3517.230 202.700 3517.370 ;
        RECT 200.200 825.870 200.460 826.190 ;
        RECT 579.700 825.870 579.960 826.190 ;
        RECT 579.760 800.000 579.900 825.870 ;
        RECT 579.490 799.270 579.900 800.000 ;
        RECT 579.490 796.000 579.770 799.270 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3416.220 17.410 3416.280 ;
        RECT 586.570 3416.220 586.890 3416.280 ;
        RECT 17.090 3416.080 586.890 3416.220 ;
        RECT 17.090 3416.020 17.410 3416.080 ;
        RECT 586.570 3416.020 586.890 3416.080 ;
      LAYER via ;
        RECT 17.120 3416.020 17.380 3416.280 ;
        RECT 586.600 3416.020 586.860 3416.280 ;
      LAYER met2 ;
        RECT 17.110 3421.235 17.390 3421.605 ;
        RECT 17.180 3416.310 17.320 3421.235 ;
        RECT 17.120 3415.990 17.380 3416.310 ;
        RECT 586.600 3415.990 586.860 3416.310 ;
        RECT 586.660 800.000 586.800 3415.990 ;
        RECT 586.390 799.270 586.800 800.000 ;
        RECT 586.390 796.000 586.670 799.270 ;
      LAYER via2 ;
        RECT 17.110 3421.280 17.390 3421.560 ;
      LAYER met3 ;
        RECT -4.800 3421.570 2.400 3422.020 ;
        RECT 17.085 3421.570 17.415 3421.585 ;
        RECT -4.800 3421.270 17.415 3421.570 ;
        RECT -4.800 3420.820 2.400 3421.270 ;
        RECT 17.085 3421.255 17.415 3421.270 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3160.540 17.410 3160.600 ;
        RECT 582.890 3160.540 583.210 3160.600 ;
        RECT 17.090 3160.400 583.210 3160.540 ;
        RECT 17.090 3160.340 17.410 3160.400 ;
        RECT 582.890 3160.340 583.210 3160.400 ;
        RECT 582.890 820.660 583.210 820.720 ;
        RECT 593.470 820.660 593.790 820.720 ;
        RECT 582.890 820.520 593.790 820.660 ;
        RECT 582.890 820.460 583.210 820.520 ;
        RECT 593.470 820.460 593.790 820.520 ;
      LAYER via ;
        RECT 17.120 3160.340 17.380 3160.600 ;
        RECT 582.920 3160.340 583.180 3160.600 ;
        RECT 582.920 820.460 583.180 820.720 ;
        RECT 593.500 820.460 593.760 820.720 ;
      LAYER met2 ;
        RECT 17.120 3160.485 17.380 3160.630 ;
        RECT 17.110 3160.115 17.390 3160.485 ;
        RECT 582.920 3160.310 583.180 3160.630 ;
        RECT 582.980 820.750 583.120 3160.310 ;
        RECT 582.920 820.430 583.180 820.750 ;
        RECT 593.500 820.430 593.760 820.750 ;
        RECT 593.560 800.000 593.700 820.430 ;
        RECT 593.290 799.270 593.700 800.000 ;
        RECT 593.290 796.000 593.570 799.270 ;
      LAYER via2 ;
        RECT 17.110 3160.160 17.390 3160.440 ;
      LAYER met3 ;
        RECT -4.800 3160.450 2.400 3160.900 ;
        RECT 17.085 3160.450 17.415 3160.465 ;
        RECT -4.800 3160.150 17.415 3160.450 ;
        RECT -4.800 3159.700 2.400 3160.150 ;
        RECT 17.085 3160.135 17.415 3160.150 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2898.400 16.950 2898.460 ;
        RECT 600.370 2898.400 600.690 2898.460 ;
        RECT 16.630 2898.260 600.690 2898.400 ;
        RECT 16.630 2898.200 16.950 2898.260 ;
        RECT 600.370 2898.200 600.690 2898.260 ;
      LAYER via ;
        RECT 16.660 2898.200 16.920 2898.460 ;
        RECT 600.400 2898.200 600.660 2898.460 ;
      LAYER met2 ;
        RECT 16.650 2899.675 16.930 2900.045 ;
        RECT 16.720 2898.490 16.860 2899.675 ;
        RECT 16.660 2898.170 16.920 2898.490 ;
        RECT 600.400 2898.170 600.660 2898.490 ;
        RECT 600.460 800.000 600.600 2898.170 ;
        RECT 600.190 799.270 600.600 800.000 ;
        RECT 600.190 796.000 600.470 799.270 ;
      LAYER via2 ;
        RECT 16.650 2899.720 16.930 2900.000 ;
      LAYER met3 ;
        RECT -4.800 2900.010 2.400 2900.460 ;
        RECT 16.625 2900.010 16.955 2900.025 ;
        RECT -4.800 2899.710 16.955 2900.010 ;
        RECT -4.800 2899.260 2.400 2899.710 ;
        RECT 16.625 2899.695 16.955 2899.710 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2635.920 17.410 2635.980 ;
        RECT 607.270 2635.920 607.590 2635.980 ;
        RECT 17.090 2635.780 607.590 2635.920 ;
        RECT 17.090 2635.720 17.410 2635.780 ;
        RECT 607.270 2635.720 607.590 2635.780 ;
      LAYER via ;
        RECT 17.120 2635.720 17.380 2635.980 ;
        RECT 607.300 2635.720 607.560 2635.980 ;
      LAYER met2 ;
        RECT 17.110 2639.235 17.390 2639.605 ;
        RECT 17.180 2636.010 17.320 2639.235 ;
        RECT 17.120 2635.690 17.380 2636.010 ;
        RECT 607.300 2635.690 607.560 2636.010 ;
        RECT 607.360 800.000 607.500 2635.690 ;
        RECT 607.090 799.270 607.500 800.000 ;
        RECT 607.090 796.000 607.370 799.270 ;
      LAYER via2 ;
        RECT 17.110 2639.280 17.390 2639.560 ;
      LAYER met3 ;
        RECT -4.800 2639.570 2.400 2640.020 ;
        RECT 17.085 2639.570 17.415 2639.585 ;
        RECT -4.800 2639.270 17.415 2639.570 ;
        RECT -4.800 2638.820 2.400 2639.270 ;
        RECT 17.085 2639.255 17.415 2639.270 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2373.780 17.410 2373.840 ;
        RECT 614.170 2373.780 614.490 2373.840 ;
        RECT 17.090 2373.640 614.490 2373.780 ;
        RECT 17.090 2373.580 17.410 2373.640 ;
        RECT 614.170 2373.580 614.490 2373.640 ;
      LAYER via ;
        RECT 17.120 2373.580 17.380 2373.840 ;
        RECT 614.200 2373.580 614.460 2373.840 ;
      LAYER met2 ;
        RECT 17.110 2378.115 17.390 2378.485 ;
        RECT 17.180 2373.870 17.320 2378.115 ;
        RECT 17.120 2373.550 17.380 2373.870 ;
        RECT 614.200 2373.550 614.460 2373.870 ;
        RECT 614.260 800.000 614.400 2373.550 ;
        RECT 613.990 799.270 614.400 800.000 ;
        RECT 613.990 796.000 614.270 799.270 ;
      LAYER via2 ;
        RECT 17.110 2378.160 17.390 2378.440 ;
      LAYER met3 ;
        RECT -4.800 2378.450 2.400 2378.900 ;
        RECT 17.085 2378.450 17.415 2378.465 ;
        RECT -4.800 2378.150 17.415 2378.450 ;
        RECT -4.800 2377.700 2.400 2378.150 ;
        RECT 17.085 2378.135 17.415 2378.150 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2111.640 17.410 2111.700 ;
        RECT 621.070 2111.640 621.390 2111.700 ;
        RECT 17.090 2111.500 621.390 2111.640 ;
        RECT 17.090 2111.440 17.410 2111.500 ;
        RECT 621.070 2111.440 621.390 2111.500 ;
      LAYER via ;
        RECT 17.120 2111.440 17.380 2111.700 ;
        RECT 621.100 2111.440 621.360 2111.700 ;
      LAYER met2 ;
        RECT 17.110 2117.675 17.390 2118.045 ;
        RECT 17.180 2111.730 17.320 2117.675 ;
        RECT 17.120 2111.410 17.380 2111.730 ;
        RECT 621.100 2111.410 621.360 2111.730 ;
        RECT 621.160 800.000 621.300 2111.410 ;
        RECT 620.890 799.270 621.300 800.000 ;
        RECT 620.890 796.000 621.170 799.270 ;
      LAYER via2 ;
        RECT 17.110 2117.720 17.390 2118.000 ;
      LAYER met3 ;
        RECT -4.800 2118.010 2.400 2118.460 ;
        RECT 17.085 2118.010 17.415 2118.025 ;
        RECT -4.800 2117.710 17.415 2118.010 ;
        RECT -4.800 2117.260 2.400 2117.710 ;
        RECT 17.085 2117.695 17.415 2117.710 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 436.150 801.280 436.470 801.340 ;
        RECT 2903.130 801.280 2903.450 801.340 ;
        RECT 436.150 801.140 2903.450 801.280 ;
        RECT 436.150 801.080 436.470 801.140 ;
        RECT 2903.130 801.080 2903.450 801.140 ;
      LAYER via ;
        RECT 436.180 801.080 436.440 801.340 ;
        RECT 2903.160 801.080 2903.420 801.340 ;
      LAYER met2 ;
        RECT 436.180 801.050 436.440 801.370 ;
        RECT 2903.160 801.050 2903.420 801.370 ;
        RECT 434.590 799.410 434.870 800.000 ;
        RECT 436.240 799.410 436.380 801.050 ;
        RECT 434.590 799.270 436.380 799.410 ;
        RECT 434.590 796.000 434.870 799.270 ;
        RECT 2903.220 430.965 2903.360 801.050 ;
        RECT 2903.150 430.595 2903.430 430.965 ;
      LAYER via2 ;
        RECT 2903.150 430.640 2903.430 430.920 ;
      LAYER met3 ;
        RECT 2903.125 430.930 2903.455 430.945 ;
        RECT 2917.600 430.930 2924.800 431.380 ;
        RECT 2903.125 430.630 2924.800 430.930 ;
        RECT 2903.125 430.615 2903.455 430.630 ;
        RECT 2917.600 430.180 2924.800 430.630 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 1856.300 17.410 1856.360 ;
        RECT 627.970 1856.300 628.290 1856.360 ;
        RECT 17.090 1856.160 628.290 1856.300 ;
        RECT 17.090 1856.100 17.410 1856.160 ;
        RECT 627.970 1856.100 628.290 1856.160 ;
      LAYER via ;
        RECT 17.120 1856.100 17.380 1856.360 ;
        RECT 628.000 1856.100 628.260 1856.360 ;
      LAYER met2 ;
        RECT 17.110 1856.555 17.390 1856.925 ;
        RECT 17.180 1856.390 17.320 1856.555 ;
        RECT 17.120 1856.070 17.380 1856.390 ;
        RECT 628.000 1856.070 628.260 1856.390 ;
        RECT 628.060 800.000 628.200 1856.070 ;
        RECT 627.790 799.270 628.200 800.000 ;
        RECT 627.790 796.000 628.070 799.270 ;
      LAYER via2 ;
        RECT 17.110 1856.600 17.390 1856.880 ;
      LAYER met3 ;
        RECT -4.800 1856.890 2.400 1857.340 ;
        RECT 17.085 1856.890 17.415 1856.905 ;
        RECT -4.800 1856.590 17.415 1856.890 ;
        RECT -4.800 1856.140 2.400 1856.590 ;
        RECT 17.085 1856.575 17.415 1856.590 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 1594.160 17.410 1594.220 ;
        RECT 634.870 1594.160 635.190 1594.220 ;
        RECT 17.090 1594.020 635.190 1594.160 ;
        RECT 17.090 1593.960 17.410 1594.020 ;
        RECT 634.870 1593.960 635.190 1594.020 ;
      LAYER via ;
        RECT 17.120 1593.960 17.380 1594.220 ;
        RECT 634.900 1593.960 635.160 1594.220 ;
      LAYER met2 ;
        RECT 17.110 1596.115 17.390 1596.485 ;
        RECT 17.180 1594.250 17.320 1596.115 ;
        RECT 17.120 1593.930 17.380 1594.250 ;
        RECT 634.900 1593.930 635.160 1594.250 ;
        RECT 634.960 800.000 635.100 1593.930 ;
        RECT 634.690 799.270 635.100 800.000 ;
        RECT 634.690 796.000 634.970 799.270 ;
      LAYER via2 ;
        RECT 17.110 1596.160 17.390 1596.440 ;
      LAYER met3 ;
        RECT -4.800 1596.450 2.400 1596.900 ;
        RECT 17.085 1596.450 17.415 1596.465 ;
        RECT -4.800 1596.150 17.415 1596.450 ;
        RECT -4.800 1595.700 2.400 1596.150 ;
        RECT 17.085 1596.135 17.415 1596.150 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 1332.020 15.570 1332.080 ;
        RECT 641.770 1332.020 642.090 1332.080 ;
        RECT 15.250 1331.880 642.090 1332.020 ;
        RECT 15.250 1331.820 15.570 1331.880 ;
        RECT 641.770 1331.820 642.090 1331.880 ;
      LAYER via ;
        RECT 15.280 1331.820 15.540 1332.080 ;
        RECT 641.800 1331.820 642.060 1332.080 ;
      LAYER met2 ;
        RECT 15.270 1335.675 15.550 1336.045 ;
        RECT 15.340 1332.110 15.480 1335.675 ;
        RECT 15.280 1331.790 15.540 1332.110 ;
        RECT 641.800 1331.790 642.060 1332.110 ;
        RECT 641.860 800.000 642.000 1331.790 ;
        RECT 641.590 799.270 642.000 800.000 ;
        RECT 641.590 796.000 641.870 799.270 ;
      LAYER via2 ;
        RECT 15.270 1335.720 15.550 1336.000 ;
      LAYER met3 ;
        RECT -4.800 1336.010 2.400 1336.460 ;
        RECT 15.245 1336.010 15.575 1336.025 ;
        RECT -4.800 1335.710 15.575 1336.010 ;
        RECT -4.800 1335.260 2.400 1335.710 ;
        RECT 15.245 1335.695 15.575 1335.710 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 1069.880 16.030 1069.940 ;
        RECT 648.670 1069.880 648.990 1069.940 ;
        RECT 15.710 1069.740 648.990 1069.880 ;
        RECT 15.710 1069.680 16.030 1069.740 ;
        RECT 648.670 1069.680 648.990 1069.740 ;
      LAYER via ;
        RECT 15.740 1069.680 16.000 1069.940 ;
        RECT 648.700 1069.680 648.960 1069.940 ;
      LAYER met2 ;
        RECT 15.730 1074.555 16.010 1074.925 ;
        RECT 15.800 1069.970 15.940 1074.555 ;
        RECT 15.740 1069.650 16.000 1069.970 ;
        RECT 648.700 1069.650 648.960 1069.970 ;
        RECT 648.760 800.000 648.900 1069.650 ;
        RECT 648.490 799.270 648.900 800.000 ;
        RECT 648.490 796.000 648.770 799.270 ;
      LAYER via2 ;
        RECT 15.730 1074.600 16.010 1074.880 ;
      LAYER met3 ;
        RECT -4.800 1074.890 2.400 1075.340 ;
        RECT 15.705 1074.890 16.035 1074.905 ;
        RECT -4.800 1074.590 16.035 1074.890 ;
        RECT -4.800 1074.140 2.400 1074.590 ;
        RECT 15.705 1074.575 16.035 1074.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 814.540 17.410 814.600 ;
        RECT 655.570 814.540 655.890 814.600 ;
        RECT 17.090 814.400 655.890 814.540 ;
        RECT 17.090 814.340 17.410 814.400 ;
        RECT 655.570 814.340 655.890 814.400 ;
      LAYER via ;
        RECT 17.120 814.340 17.380 814.600 ;
        RECT 655.600 814.340 655.860 814.600 ;
      LAYER met2 ;
        RECT 17.120 814.485 17.380 814.630 ;
        RECT 17.110 814.115 17.390 814.485 ;
        RECT 655.600 814.310 655.860 814.630 ;
        RECT 655.660 800.000 655.800 814.310 ;
        RECT 655.390 799.270 655.800 800.000 ;
        RECT 655.390 796.000 655.670 799.270 ;
      LAYER via2 ;
        RECT 17.110 814.160 17.390 814.440 ;
      LAYER met3 ;
        RECT -4.800 814.450 2.400 814.900 ;
        RECT 17.085 814.450 17.415 814.465 ;
        RECT -4.800 814.150 17.415 814.450 ;
        RECT -4.800 813.700 2.400 814.150 ;
        RECT 17.085 814.135 17.415 814.150 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.930 802.980 19.250 803.040 ;
        RECT 662.470 802.980 662.790 803.040 ;
        RECT 18.930 802.840 662.790 802.980 ;
        RECT 18.930 802.780 19.250 802.840 ;
        RECT 662.470 802.780 662.790 802.840 ;
      LAYER via ;
        RECT 18.960 802.780 19.220 803.040 ;
        RECT 662.500 802.780 662.760 803.040 ;
      LAYER met2 ;
        RECT 18.960 802.750 19.220 803.070 ;
        RECT 662.500 802.750 662.760 803.070 ;
        RECT 19.020 553.365 19.160 802.750 ;
        RECT 662.560 800.000 662.700 802.750 ;
        RECT 662.290 799.270 662.700 800.000 ;
        RECT 662.290 796.000 662.570 799.270 ;
        RECT 18.950 552.995 19.230 553.365 ;
      LAYER via2 ;
        RECT 18.950 553.040 19.230 553.320 ;
      LAYER met3 ;
        RECT -4.800 553.330 2.400 553.780 ;
        RECT 18.925 553.330 19.255 553.345 ;
        RECT -4.800 553.030 19.255 553.330 ;
        RECT -4.800 552.580 2.400 553.030 ;
        RECT 18.925 553.015 19.255 553.030 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.470 802.640 18.790 802.700 ;
        RECT 669.370 802.640 669.690 802.700 ;
        RECT 18.470 802.500 669.690 802.640 ;
        RECT 18.470 802.440 18.790 802.500 ;
        RECT 669.370 802.440 669.690 802.500 ;
      LAYER via ;
        RECT 18.500 802.440 18.760 802.700 ;
        RECT 669.400 802.440 669.660 802.700 ;
      LAYER met2 ;
        RECT 18.500 802.410 18.760 802.730 ;
        RECT 669.400 802.410 669.660 802.730 ;
        RECT 18.560 358.205 18.700 802.410 ;
        RECT 669.460 800.000 669.600 802.410 ;
        RECT 669.190 799.270 669.600 800.000 ;
        RECT 669.190 796.000 669.470 799.270 ;
        RECT 18.490 357.835 18.770 358.205 ;
      LAYER via2 ;
        RECT 18.490 357.880 18.770 358.160 ;
      LAYER met3 ;
        RECT -4.800 358.170 2.400 358.620 ;
        RECT 18.465 358.170 18.795 358.185 ;
        RECT -4.800 357.870 18.795 358.170 ;
        RECT -4.800 357.420 2.400 357.870 ;
        RECT 18.465 357.855 18.795 357.870 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 801.960 17.410 802.020 ;
        RECT 676.270 801.960 676.590 802.020 ;
        RECT 17.090 801.820 676.590 801.960 ;
        RECT 17.090 801.760 17.410 801.820 ;
        RECT 676.270 801.760 676.590 801.820 ;
      LAYER via ;
        RECT 17.120 801.760 17.380 802.020 ;
        RECT 676.300 801.760 676.560 802.020 ;
      LAYER met2 ;
        RECT 17.120 801.730 17.380 802.050 ;
        RECT 676.300 801.730 676.560 802.050 ;
        RECT 17.180 162.365 17.320 801.730 ;
        RECT 676.360 800.000 676.500 801.730 ;
        RECT 676.090 799.270 676.500 800.000 ;
        RECT 676.090 796.000 676.370 799.270 ;
        RECT 17.110 161.995 17.390 162.365 ;
      LAYER via2 ;
        RECT 17.110 162.040 17.390 162.320 ;
      LAYER met3 ;
        RECT -4.800 162.330 2.400 162.780 ;
        RECT 17.085 162.330 17.415 162.345 ;
        RECT -4.800 162.030 17.415 162.330 ;
        RECT -4.800 161.580 2.400 162.030 ;
        RECT 17.085 162.015 17.415 162.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 443.050 801.620 443.370 801.680 ;
        RECT 2904.050 801.620 2904.370 801.680 ;
        RECT 443.050 801.480 2904.370 801.620 ;
        RECT 443.050 801.420 443.370 801.480 ;
        RECT 2904.050 801.420 2904.370 801.480 ;
      LAYER via ;
        RECT 443.080 801.420 443.340 801.680 ;
        RECT 2904.080 801.420 2904.340 801.680 ;
      LAYER met2 ;
        RECT 443.080 801.390 443.340 801.710 ;
        RECT 2904.080 801.390 2904.340 801.710 ;
        RECT 441.490 799.410 441.770 800.000 ;
        RECT 443.140 799.410 443.280 801.390 ;
        RECT 441.490 799.270 443.280 799.410 ;
        RECT 441.490 796.000 441.770 799.270 ;
        RECT 2904.140 630.205 2904.280 801.390 ;
        RECT 2904.070 629.835 2904.350 630.205 ;
      LAYER via2 ;
        RECT 2904.070 629.880 2904.350 630.160 ;
      LAYER met3 ;
        RECT 2904.045 630.170 2904.375 630.185 ;
        RECT 2917.600 630.170 2924.800 630.620 ;
        RECT 2904.045 629.870 2924.800 630.170 ;
        RECT 2904.045 629.855 2904.375 629.870 ;
        RECT 2917.600 629.420 2924.800 629.870 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.570 828.140 448.890 828.200 ;
        RECT 2900.830 828.140 2901.150 828.200 ;
        RECT 448.570 828.000 2901.150 828.140 ;
        RECT 448.570 827.940 448.890 828.000 ;
        RECT 2900.830 827.940 2901.150 828.000 ;
      LAYER via ;
        RECT 448.600 827.940 448.860 828.200 ;
        RECT 2900.860 827.940 2901.120 828.200 ;
      LAYER met2 ;
        RECT 2900.850 829.075 2901.130 829.445 ;
        RECT 2900.920 828.230 2901.060 829.075 ;
        RECT 448.600 827.910 448.860 828.230 ;
        RECT 2900.860 827.910 2901.120 828.230 ;
        RECT 448.660 800.000 448.800 827.910 ;
        RECT 448.390 799.270 448.800 800.000 ;
        RECT 448.390 796.000 448.670 799.270 ;
      LAYER via2 ;
        RECT 2900.850 829.120 2901.130 829.400 ;
      LAYER met3 ;
        RECT 2900.825 829.410 2901.155 829.425 ;
        RECT 2917.600 829.410 2924.800 829.860 ;
        RECT 2900.825 829.110 2924.800 829.410 ;
        RECT 2900.825 829.095 2901.155 829.110 ;
        RECT 2917.600 828.660 2924.800 829.110 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.470 1028.400 455.790 1028.460 ;
        RECT 2900.830 1028.400 2901.150 1028.460 ;
        RECT 455.470 1028.260 2901.150 1028.400 ;
        RECT 455.470 1028.200 455.790 1028.260 ;
        RECT 2900.830 1028.200 2901.150 1028.260 ;
      LAYER via ;
        RECT 455.500 1028.200 455.760 1028.460 ;
        RECT 2900.860 1028.200 2901.120 1028.460 ;
      LAYER met2 ;
        RECT 455.500 1028.170 455.760 1028.490 ;
        RECT 2900.850 1028.315 2901.130 1028.685 ;
        RECT 2900.860 1028.170 2901.120 1028.315 ;
        RECT 455.560 800.000 455.700 1028.170 ;
        RECT 455.290 799.270 455.700 800.000 ;
        RECT 455.290 796.000 455.570 799.270 ;
      LAYER via2 ;
        RECT 2900.850 1028.360 2901.130 1028.640 ;
      LAYER met3 ;
        RECT 2900.825 1028.650 2901.155 1028.665 ;
        RECT 2917.600 1028.650 2924.800 1029.100 ;
        RECT 2900.825 1028.350 2924.800 1028.650 ;
        RECT 2900.825 1028.335 2901.155 1028.350 ;
        RECT 2917.600 1027.900 2924.800 1028.350 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.370 1221.520 462.690 1221.580 ;
        RECT 2898.990 1221.520 2899.310 1221.580 ;
        RECT 462.370 1221.380 2899.310 1221.520 ;
        RECT 462.370 1221.320 462.690 1221.380 ;
        RECT 2898.990 1221.320 2899.310 1221.380 ;
      LAYER via ;
        RECT 462.400 1221.320 462.660 1221.580 ;
        RECT 2899.020 1221.320 2899.280 1221.580 ;
      LAYER met2 ;
        RECT 2899.010 1227.555 2899.290 1227.925 ;
        RECT 2899.080 1221.610 2899.220 1227.555 ;
        RECT 462.400 1221.290 462.660 1221.610 ;
        RECT 2899.020 1221.290 2899.280 1221.610 ;
        RECT 462.460 800.000 462.600 1221.290 ;
        RECT 462.190 799.270 462.600 800.000 ;
        RECT 462.190 796.000 462.470 799.270 ;
      LAYER via2 ;
        RECT 2899.010 1227.600 2899.290 1227.880 ;
      LAYER met3 ;
        RECT 2898.985 1227.890 2899.315 1227.905 ;
        RECT 2917.600 1227.890 2924.800 1228.340 ;
        RECT 2898.985 1227.590 2924.800 1227.890 ;
        RECT 2898.985 1227.575 2899.315 1227.590 ;
        RECT 2917.600 1227.140 2924.800 1227.590 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.270 1490.800 469.590 1490.860 ;
        RECT 2900.830 1490.800 2901.150 1490.860 ;
        RECT 469.270 1490.660 2901.150 1490.800 ;
        RECT 469.270 1490.600 469.590 1490.660 ;
        RECT 2900.830 1490.600 2901.150 1490.660 ;
      LAYER via ;
        RECT 469.300 1490.600 469.560 1490.860 ;
        RECT 2900.860 1490.600 2901.120 1490.860 ;
      LAYER met2 ;
        RECT 2900.850 1493.435 2901.130 1493.805 ;
        RECT 2900.920 1490.890 2901.060 1493.435 ;
        RECT 469.300 1490.570 469.560 1490.890 ;
        RECT 2900.860 1490.570 2901.120 1490.890 ;
        RECT 469.360 800.000 469.500 1490.570 ;
        RECT 469.090 799.270 469.500 800.000 ;
        RECT 469.090 796.000 469.370 799.270 ;
      LAYER via2 ;
        RECT 2900.850 1493.480 2901.130 1493.760 ;
      LAYER met3 ;
        RECT 2900.825 1493.770 2901.155 1493.785 ;
        RECT 2917.600 1493.770 2924.800 1494.220 ;
        RECT 2900.825 1493.470 2924.800 1493.770 ;
        RECT 2900.825 1493.455 2901.155 1493.470 ;
        RECT 2917.600 1493.020 2924.800 1493.470 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.170 1759.740 476.490 1759.800 ;
        RECT 2900.830 1759.740 2901.150 1759.800 ;
        RECT 476.170 1759.600 2901.150 1759.740 ;
        RECT 476.170 1759.540 476.490 1759.600 ;
        RECT 2900.830 1759.540 2901.150 1759.600 ;
      LAYER via ;
        RECT 476.200 1759.540 476.460 1759.800 ;
        RECT 2900.860 1759.540 2901.120 1759.800 ;
      LAYER met2 ;
        RECT 476.200 1759.510 476.460 1759.830 ;
        RECT 2900.860 1759.685 2901.120 1759.830 ;
        RECT 476.260 800.000 476.400 1759.510 ;
        RECT 2900.850 1759.315 2901.130 1759.685 ;
        RECT 475.990 799.270 476.400 800.000 ;
        RECT 475.990 796.000 476.270 799.270 ;
      LAYER via2 ;
        RECT 2900.850 1759.360 2901.130 1759.640 ;
      LAYER met3 ;
        RECT 2900.825 1759.650 2901.155 1759.665 ;
        RECT 2917.600 1759.650 2924.800 1760.100 ;
        RECT 2900.825 1759.350 2924.800 1759.650 ;
        RECT 2900.825 1759.335 2901.155 1759.350 ;
        RECT 2917.600 1758.900 2924.800 1759.350 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.070 2021.880 483.390 2021.940 ;
        RECT 2900.830 2021.880 2901.150 2021.940 ;
        RECT 483.070 2021.740 2901.150 2021.880 ;
        RECT 483.070 2021.680 483.390 2021.740 ;
        RECT 2900.830 2021.680 2901.150 2021.740 ;
      LAYER via ;
        RECT 483.100 2021.680 483.360 2021.940 ;
        RECT 2900.860 2021.680 2901.120 2021.940 ;
      LAYER met2 ;
        RECT 2900.850 2024.515 2901.130 2024.885 ;
        RECT 2900.920 2021.970 2901.060 2024.515 ;
        RECT 483.100 2021.650 483.360 2021.970 ;
        RECT 2900.860 2021.650 2901.120 2021.970 ;
        RECT 483.160 800.000 483.300 2021.650 ;
        RECT 482.890 799.270 483.300 800.000 ;
        RECT 482.890 796.000 483.170 799.270 ;
      LAYER via2 ;
        RECT 2900.850 2024.560 2901.130 2024.840 ;
      LAYER met3 ;
        RECT 2900.825 2024.850 2901.155 2024.865 ;
        RECT 2917.600 2024.850 2924.800 2025.300 ;
        RECT 2900.825 2024.550 2924.800 2024.850 ;
        RECT 2900.825 2024.535 2901.155 2024.550 ;
        RECT 2917.600 2024.100 2924.800 2024.550 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 424.190 796.660 424.510 796.920 ;
        RECT 424.280 793.460 424.420 796.660 ;
        RECT 2901.750 793.800 2902.070 793.860 ;
        RECT 469.130 793.660 2902.070 793.800 ;
        RECT 469.130 793.460 469.270 793.660 ;
        RECT 2901.750 793.600 2902.070 793.660 ;
        RECT 424.280 793.320 469.270 793.460 ;
      LAYER via ;
        RECT 424.220 796.660 424.480 796.920 ;
        RECT 2901.780 793.600 2902.040 793.860 ;
      LAYER met2 ;
        RECT 423.090 796.690 423.370 800.000 ;
        RECT 424.220 796.690 424.480 796.950 ;
        RECT 423.090 796.630 424.480 796.690 ;
        RECT 423.090 796.550 424.420 796.630 ;
        RECT 423.090 796.000 423.370 796.550 ;
        RECT 2901.780 793.570 2902.040 793.890 ;
        RECT 2901.840 165.765 2901.980 793.570 ;
        RECT 2901.770 165.395 2902.050 165.765 ;
      LAYER via2 ;
        RECT 2901.770 165.440 2902.050 165.720 ;
      LAYER met3 ;
        RECT 2901.745 165.730 2902.075 165.745 ;
        RECT 2917.600 165.730 2924.800 166.180 ;
        RECT 2901.745 165.430 2924.800 165.730 ;
        RECT 2901.745 165.415 2902.075 165.430 ;
        RECT 2917.600 164.980 2924.800 165.430 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.430 2422.060 490.750 2422.120 ;
        RECT 2900.830 2422.060 2901.150 2422.120 ;
        RECT 490.430 2421.920 2901.150 2422.060 ;
        RECT 490.430 2421.860 490.750 2421.920 ;
        RECT 2900.830 2421.860 2901.150 2421.920 ;
      LAYER via ;
        RECT 490.460 2421.860 490.720 2422.120 ;
        RECT 2900.860 2421.860 2901.120 2422.120 ;
      LAYER met2 ;
        RECT 2900.850 2422.995 2901.130 2423.365 ;
        RECT 2900.920 2422.150 2901.060 2422.995 ;
        RECT 490.460 2421.830 490.720 2422.150 ;
        RECT 2900.860 2421.830 2901.120 2422.150 ;
        RECT 490.520 799.410 490.660 2421.830 ;
        RECT 492.090 799.410 492.370 800.000 ;
        RECT 490.520 799.270 492.370 799.410 ;
        RECT 492.090 796.000 492.370 799.270 ;
      LAYER via2 ;
        RECT 2900.850 2423.040 2901.130 2423.320 ;
      LAYER met3 ;
        RECT 2900.825 2423.330 2901.155 2423.345 ;
        RECT 2917.600 2423.330 2924.800 2423.780 ;
        RECT 2900.825 2423.030 2924.800 2423.330 ;
        RECT 2900.825 2423.015 2901.155 2423.030 ;
        RECT 2917.600 2422.580 2924.800 2423.030 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.330 2684.200 497.650 2684.260 ;
        RECT 2900.830 2684.200 2901.150 2684.260 ;
        RECT 497.330 2684.060 2901.150 2684.200 ;
        RECT 497.330 2684.000 497.650 2684.060 ;
        RECT 2900.830 2684.000 2901.150 2684.060 ;
      LAYER via ;
        RECT 497.360 2684.000 497.620 2684.260 ;
        RECT 2900.860 2684.000 2901.120 2684.260 ;
      LAYER met2 ;
        RECT 2900.850 2688.875 2901.130 2689.245 ;
        RECT 2900.920 2684.290 2901.060 2688.875 ;
        RECT 497.360 2683.970 497.620 2684.290 ;
        RECT 2900.860 2683.970 2901.120 2684.290 ;
        RECT 497.420 799.410 497.560 2683.970 ;
        RECT 498.990 799.410 499.270 800.000 ;
        RECT 497.420 799.270 499.270 799.410 ;
        RECT 498.990 796.000 499.270 799.270 ;
      LAYER via2 ;
        RECT 2900.850 2688.920 2901.130 2689.200 ;
      LAYER met3 ;
        RECT 2900.825 2689.210 2901.155 2689.225 ;
        RECT 2917.600 2689.210 2924.800 2689.660 ;
        RECT 2900.825 2688.910 2924.800 2689.210 ;
        RECT 2900.825 2688.895 2901.155 2688.910 ;
        RECT 2917.600 2688.460 2924.800 2688.910 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.230 2953.480 504.550 2953.540 ;
        RECT 2898.990 2953.480 2899.310 2953.540 ;
        RECT 504.230 2953.340 2899.310 2953.480 ;
        RECT 504.230 2953.280 504.550 2953.340 ;
        RECT 2898.990 2953.280 2899.310 2953.340 ;
      LAYER via ;
        RECT 504.260 2953.280 504.520 2953.540 ;
        RECT 2899.020 2953.280 2899.280 2953.540 ;
      LAYER met2 ;
        RECT 2899.010 2954.755 2899.290 2955.125 ;
        RECT 2899.080 2953.570 2899.220 2954.755 ;
        RECT 504.260 2953.250 504.520 2953.570 ;
        RECT 2899.020 2953.250 2899.280 2953.570 ;
        RECT 504.320 799.410 504.460 2953.250 ;
        RECT 505.890 799.410 506.170 800.000 ;
        RECT 504.320 799.270 506.170 799.410 ;
        RECT 505.890 796.000 506.170 799.270 ;
      LAYER via2 ;
        RECT 2899.010 2954.800 2899.290 2955.080 ;
      LAYER met3 ;
        RECT 2898.985 2955.090 2899.315 2955.105 ;
        RECT 2917.600 2955.090 2924.800 2955.540 ;
        RECT 2898.985 2954.790 2924.800 2955.090 ;
        RECT 2898.985 2954.775 2899.315 2954.790 ;
        RECT 2917.600 2954.340 2924.800 2954.790 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.130 3215.620 511.450 3215.680 ;
        RECT 2900.830 3215.620 2901.150 3215.680 ;
        RECT 511.130 3215.480 2901.150 3215.620 ;
        RECT 511.130 3215.420 511.450 3215.480 ;
        RECT 2900.830 3215.420 2901.150 3215.480 ;
      LAYER via ;
        RECT 511.160 3215.420 511.420 3215.680 ;
        RECT 2900.860 3215.420 2901.120 3215.680 ;
      LAYER met2 ;
        RECT 2900.850 3219.955 2901.130 3220.325 ;
        RECT 2900.920 3215.710 2901.060 3219.955 ;
        RECT 511.160 3215.390 511.420 3215.710 ;
        RECT 2900.860 3215.390 2901.120 3215.710 ;
        RECT 511.220 799.410 511.360 3215.390 ;
        RECT 512.790 799.410 513.070 800.000 ;
        RECT 511.220 799.270 513.070 799.410 ;
        RECT 512.790 796.000 513.070 799.270 ;
      LAYER via2 ;
        RECT 2900.850 3220.000 2901.130 3220.280 ;
      LAYER met3 ;
        RECT 2900.825 3220.290 2901.155 3220.305 ;
        RECT 2917.600 3220.290 2924.800 3220.740 ;
        RECT 2900.825 3219.990 2924.800 3220.290 ;
        RECT 2900.825 3219.975 2901.155 3219.990 ;
        RECT 2917.600 3219.540 2924.800 3219.990 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.030 3484.900 518.350 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 518.030 3484.760 2901.150 3484.900 ;
        RECT 518.030 3484.700 518.350 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 518.060 3484.700 518.320 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3485.835 2901.130 3486.205 ;
        RECT 2900.920 3484.990 2901.060 3485.835 ;
        RECT 518.060 3484.670 518.320 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 518.120 799.410 518.260 3484.670 ;
        RECT 519.690 799.410 519.970 800.000 ;
        RECT 518.120 799.270 519.970 799.410 ;
        RECT 519.690 796.000 519.970 799.270 ;
      LAYER via2 ;
        RECT 2900.850 3485.880 2901.130 3486.160 ;
      LAYER met3 ;
        RECT 2900.825 3486.170 2901.155 3486.185 ;
        RECT 2917.600 3486.170 2924.800 3486.620 ;
        RECT 2900.825 3485.870 2924.800 3486.170 ;
        RECT 2900.825 3485.855 2901.155 3485.870 ;
        RECT 2917.600 3485.420 2924.800 3485.870 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.930 824.400 525.250 824.460 ;
        RECT 2635.870 824.400 2636.190 824.460 ;
        RECT 524.930 824.260 2636.190 824.400 ;
        RECT 524.930 824.200 525.250 824.260 ;
        RECT 2635.870 824.200 2636.190 824.260 ;
      LAYER via ;
        RECT 524.960 824.200 525.220 824.460 ;
        RECT 2635.900 824.200 2636.160 824.460 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 824.490 2636.100 3517.600 ;
        RECT 524.960 824.170 525.220 824.490 ;
        RECT 2635.900 824.170 2636.160 824.490 ;
        RECT 525.020 799.410 525.160 824.170 ;
        RECT 526.590 799.410 526.870 800.000 ;
        RECT 525.020 799.270 526.870 799.410 ;
        RECT 526.590 796.000 526.870 799.270 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 532.290 824.740 532.610 824.800 ;
        RECT 2311.570 824.740 2311.890 824.800 ;
        RECT 532.290 824.600 2311.890 824.740 ;
        RECT 532.290 824.540 532.610 824.600 ;
        RECT 2311.570 824.540 2311.890 824.600 ;
      LAYER via ;
        RECT 532.320 824.540 532.580 824.800 ;
        RECT 2311.600 824.540 2311.860 824.800 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 824.830 2311.800 3517.600 ;
        RECT 532.320 824.510 532.580 824.830 ;
        RECT 2311.600 824.510 2311.860 824.830 ;
        RECT 532.380 799.410 532.520 824.510 ;
        RECT 533.490 799.410 533.770 800.000 ;
        RECT 532.380 799.270 533.770 799.410 ;
        RECT 533.490 796.000 533.770 799.270 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 539.190 825.080 539.510 825.140 ;
        RECT 1987.270 825.080 1987.590 825.140 ;
        RECT 539.190 824.940 1987.590 825.080 ;
        RECT 539.190 824.880 539.510 824.940 ;
        RECT 1987.270 824.880 1987.590 824.940 ;
      LAYER via ;
        RECT 539.220 824.880 539.480 825.140 ;
        RECT 1987.300 824.880 1987.560 825.140 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 825.170 1987.500 3517.600 ;
        RECT 539.220 824.850 539.480 825.170 ;
        RECT 1987.300 824.850 1987.560 825.170 ;
        RECT 539.280 799.410 539.420 824.850 ;
        RECT 540.390 799.410 540.670 800.000 ;
        RECT 539.280 799.270 540.670 799.410 ;
        RECT 540.390 796.000 540.670 799.270 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1656.070 3515.160 1656.390 3515.220 ;
        RECT 1662.510 3515.160 1662.830 3515.220 ;
        RECT 1656.070 3515.020 1662.830 3515.160 ;
        RECT 1656.070 3514.960 1656.390 3515.020 ;
        RECT 1662.510 3514.960 1662.830 3515.020 ;
        RECT 545.630 825.420 545.950 825.480 ;
        RECT 1656.070 825.420 1656.390 825.480 ;
        RECT 545.630 825.280 1656.390 825.420 ;
        RECT 545.630 825.220 545.950 825.280 ;
        RECT 1656.070 825.220 1656.390 825.280 ;
      LAYER via ;
        RECT 1656.100 3514.960 1656.360 3515.220 ;
        RECT 1662.540 3514.960 1662.800 3515.220 ;
        RECT 545.660 825.220 545.920 825.480 ;
        RECT 1656.100 825.220 1656.360 825.480 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3515.250 1662.740 3517.600 ;
        RECT 1656.100 3514.930 1656.360 3515.250 ;
        RECT 1662.540 3514.930 1662.800 3515.250 ;
        RECT 1656.160 825.510 1656.300 3514.930 ;
        RECT 545.660 825.190 545.920 825.510 ;
        RECT 1656.100 825.190 1656.360 825.510 ;
        RECT 545.720 799.410 545.860 825.190 ;
        RECT 547.290 799.410 547.570 800.000 ;
        RECT 545.720 799.270 547.570 799.410 ;
        RECT 547.290 796.000 547.570 799.270 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1331.770 3487.960 1332.090 3488.020 ;
        RECT 1338.210 3487.960 1338.530 3488.020 ;
        RECT 1331.770 3487.820 1338.530 3487.960 ;
        RECT 1331.770 3487.760 1332.090 3487.820 ;
        RECT 1338.210 3487.760 1338.530 3487.820 ;
        RECT 552.990 825.760 553.310 825.820 ;
        RECT 1331.770 825.760 1332.090 825.820 ;
        RECT 552.990 825.620 1332.090 825.760 ;
        RECT 552.990 825.560 553.310 825.620 ;
        RECT 1331.770 825.560 1332.090 825.620 ;
      LAYER via ;
        RECT 1331.800 3487.760 1332.060 3488.020 ;
        RECT 1338.240 3487.760 1338.500 3488.020 ;
        RECT 553.020 825.560 553.280 825.820 ;
        RECT 1331.800 825.560 1332.060 825.820 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3488.050 1338.440 3517.600 ;
        RECT 1331.800 3487.730 1332.060 3488.050 ;
        RECT 1338.240 3487.730 1338.500 3488.050 ;
        RECT 1331.860 825.850 1332.000 3487.730 ;
        RECT 553.020 825.530 553.280 825.850 ;
        RECT 1331.800 825.530 1332.060 825.850 ;
        RECT 553.080 799.410 553.220 825.530 ;
        RECT 554.190 799.410 554.470 800.000 ;
        RECT 553.080 799.270 554.470 799.410 ;
        RECT 554.190 796.000 554.470 799.270 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 431.550 803.320 431.870 803.380 ;
        RECT 686.390 803.320 686.710 803.380 ;
        RECT 431.550 803.180 686.710 803.320 ;
        RECT 431.550 803.120 431.870 803.180 ;
        RECT 686.390 803.120 686.710 803.180 ;
        RECT 686.390 365.740 686.710 365.800 ;
        RECT 2898.070 365.740 2898.390 365.800 ;
        RECT 686.390 365.600 2898.390 365.740 ;
        RECT 686.390 365.540 686.710 365.600 ;
        RECT 2898.070 365.540 2898.390 365.600 ;
      LAYER via ;
        RECT 431.580 803.120 431.840 803.380 ;
        RECT 686.420 803.120 686.680 803.380 ;
        RECT 686.420 365.540 686.680 365.800 ;
        RECT 2898.100 365.540 2898.360 365.800 ;
      LAYER met2 ;
        RECT 431.580 803.090 431.840 803.410 ;
        RECT 686.420 803.090 686.680 803.410 ;
        RECT 429.990 799.410 430.270 800.000 ;
        RECT 431.640 799.410 431.780 803.090 ;
        RECT 429.990 799.270 431.780 799.410 ;
        RECT 429.990 796.000 430.270 799.270 ;
        RECT 686.480 365.830 686.620 803.090 ;
        RECT 686.420 365.510 686.680 365.830 ;
        RECT 2898.100 365.510 2898.360 365.830 ;
        RECT 2898.160 365.005 2898.300 365.510 ;
        RECT 2898.090 364.635 2898.370 365.005 ;
      LAYER via2 ;
        RECT 2898.090 364.680 2898.370 364.960 ;
      LAYER met3 ;
        RECT 2898.065 364.970 2898.395 364.985 ;
        RECT 2917.600 364.970 2924.800 365.420 ;
        RECT 2898.065 364.670 2924.800 364.970 ;
        RECT 2898.065 364.655 2898.395 364.670 ;
        RECT 2917.600 364.220 2924.800 364.670 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.430 3502.920 559.750 3502.980 ;
        RECT 1013.910 3502.920 1014.230 3502.980 ;
        RECT 559.430 3502.780 1014.230 3502.920 ;
        RECT 559.430 3502.720 559.750 3502.780 ;
        RECT 1013.910 3502.720 1014.230 3502.780 ;
      LAYER via ;
        RECT 559.460 3502.720 559.720 3502.980 ;
        RECT 1013.940 3502.720 1014.200 3502.980 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3503.010 1014.140 3517.600 ;
        RECT 559.460 3502.690 559.720 3503.010 ;
        RECT 1013.940 3502.690 1014.200 3503.010 ;
        RECT 559.520 799.410 559.660 3502.690 ;
        RECT 561.090 799.410 561.370 800.000 ;
        RECT 559.520 799.270 561.370 799.410 ;
        RECT 561.090 796.000 561.370 799.270 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.330 3503.260 566.650 3503.320 ;
        RECT 689.150 3503.260 689.470 3503.320 ;
        RECT 566.330 3503.120 689.470 3503.260 ;
        RECT 566.330 3503.060 566.650 3503.120 ;
        RECT 689.150 3503.060 689.470 3503.120 ;
      LAYER via ;
        RECT 566.360 3503.060 566.620 3503.320 ;
        RECT 689.180 3503.060 689.440 3503.320 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3503.350 689.380 3517.600 ;
        RECT 566.360 3503.030 566.620 3503.350 ;
        RECT 689.180 3503.030 689.440 3503.350 ;
        RECT 566.420 799.410 566.560 3503.030 ;
        RECT 567.990 799.410 568.270 800.000 ;
        RECT 566.420 799.270 568.270 799.410 ;
        RECT 567.990 796.000 568.270 799.270 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 358.870 3515.160 359.190 3515.220 ;
        RECT 364.850 3515.160 365.170 3515.220 ;
        RECT 358.870 3515.020 365.170 3515.160 ;
        RECT 358.870 3514.960 359.190 3515.020 ;
        RECT 364.850 3514.960 365.170 3515.020 ;
        RECT 358.870 826.780 359.190 826.840 ;
        RECT 573.230 826.780 573.550 826.840 ;
        RECT 358.870 826.640 573.550 826.780 ;
        RECT 358.870 826.580 359.190 826.640 ;
        RECT 573.230 826.580 573.550 826.640 ;
      LAYER via ;
        RECT 358.900 3514.960 359.160 3515.220 ;
        RECT 364.880 3514.960 365.140 3515.220 ;
        RECT 358.900 826.580 359.160 826.840 ;
        RECT 573.260 826.580 573.520 826.840 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3515.250 365.080 3517.600 ;
        RECT 358.900 3514.930 359.160 3515.250 ;
        RECT 364.880 3514.930 365.140 3515.250 ;
        RECT 358.960 826.870 359.100 3514.930 ;
        RECT 358.900 826.550 359.160 826.870 ;
        RECT 573.260 826.550 573.520 826.870 ;
        RECT 573.320 799.410 573.460 826.550 ;
        RECT 574.890 799.410 575.170 800.000 ;
        RECT 573.320 799.270 575.170 799.410 ;
        RECT 574.890 796.000 575.170 799.270 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.570 831.880 34.890 831.940 ;
        RECT 580.130 831.880 580.450 831.940 ;
        RECT 34.570 831.740 580.450 831.880 ;
        RECT 34.570 831.680 34.890 831.740 ;
        RECT 580.130 831.680 580.450 831.740 ;
      LAYER via ;
        RECT 34.600 831.680 34.860 831.940 ;
        RECT 580.160 831.680 580.420 831.940 ;
      LAYER met2 ;
        RECT 34.660 3517.910 39.860 3518.050 ;
        RECT 34.660 831.970 34.800 3517.910 ;
        RECT 39.720 3517.370 39.860 3517.910 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3517.370 40.780 3517.600 ;
        RECT 39.720 3517.230 40.780 3517.370 ;
        RECT 34.600 831.650 34.860 831.970 ;
        RECT 580.160 831.650 580.420 831.970 ;
        RECT 580.220 799.410 580.360 831.650 ;
        RECT 581.790 799.410 582.070 800.000 ;
        RECT 580.220 799.270 582.070 799.410 ;
        RECT 581.790 796.000 582.070 799.270 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3284.640 17.410 3284.700 ;
        RECT 587.490 3284.640 587.810 3284.700 ;
        RECT 17.090 3284.500 587.810 3284.640 ;
        RECT 17.090 3284.440 17.410 3284.500 ;
        RECT 587.490 3284.440 587.810 3284.500 ;
      LAYER via ;
        RECT 17.120 3284.440 17.380 3284.700 ;
        RECT 587.520 3284.440 587.780 3284.700 ;
      LAYER met2 ;
        RECT 17.110 3290.675 17.390 3291.045 ;
        RECT 17.180 3284.730 17.320 3290.675 ;
        RECT 17.120 3284.410 17.380 3284.730 ;
        RECT 587.520 3284.410 587.780 3284.730 ;
        RECT 587.580 799.410 587.720 3284.410 ;
        RECT 588.690 799.410 588.970 800.000 ;
        RECT 587.580 799.270 588.970 799.410 ;
        RECT 588.690 796.000 588.970 799.270 ;
      LAYER via2 ;
        RECT 17.110 3290.720 17.390 3291.000 ;
      LAYER met3 ;
        RECT -4.800 3291.010 2.400 3291.460 ;
        RECT 17.085 3291.010 17.415 3291.025 ;
        RECT -4.800 3290.710 17.415 3291.010 ;
        RECT -4.800 3290.260 2.400 3290.710 ;
        RECT 17.085 3290.695 17.415 3290.710 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 3029.300 16.490 3029.360 ;
        RECT 594.390 3029.300 594.710 3029.360 ;
        RECT 16.170 3029.160 594.710 3029.300 ;
        RECT 16.170 3029.100 16.490 3029.160 ;
        RECT 594.390 3029.100 594.710 3029.160 ;
      LAYER via ;
        RECT 16.200 3029.100 16.460 3029.360 ;
        RECT 594.420 3029.100 594.680 3029.360 ;
      LAYER met2 ;
        RECT 16.190 3030.235 16.470 3030.605 ;
        RECT 16.260 3029.390 16.400 3030.235 ;
        RECT 16.200 3029.070 16.460 3029.390 ;
        RECT 594.420 3029.070 594.680 3029.390 ;
        RECT 594.480 799.410 594.620 3029.070 ;
        RECT 595.590 799.410 595.870 800.000 ;
        RECT 594.480 799.270 595.870 799.410 ;
        RECT 595.590 796.000 595.870 799.270 ;
      LAYER via2 ;
        RECT 16.190 3030.280 16.470 3030.560 ;
      LAYER met3 ;
        RECT -4.800 3030.570 2.400 3031.020 ;
        RECT 16.165 3030.570 16.495 3030.585 ;
        RECT -4.800 3030.270 16.495 3030.570 ;
        RECT -4.800 3029.820 2.400 3030.270 ;
        RECT 16.165 3030.255 16.495 3030.270 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2767.160 17.410 2767.220 ;
        RECT 601.290 2767.160 601.610 2767.220 ;
        RECT 17.090 2767.020 601.610 2767.160 ;
        RECT 17.090 2766.960 17.410 2767.020 ;
        RECT 601.290 2766.960 601.610 2767.020 ;
      LAYER via ;
        RECT 17.120 2766.960 17.380 2767.220 ;
        RECT 601.320 2766.960 601.580 2767.220 ;
      LAYER met2 ;
        RECT 17.110 2769.115 17.390 2769.485 ;
        RECT 17.180 2767.250 17.320 2769.115 ;
        RECT 17.120 2766.930 17.380 2767.250 ;
        RECT 601.320 2766.930 601.580 2767.250 ;
        RECT 601.380 799.410 601.520 2766.930 ;
        RECT 602.490 799.410 602.770 800.000 ;
        RECT 601.380 799.270 602.770 799.410 ;
        RECT 602.490 796.000 602.770 799.270 ;
      LAYER via2 ;
        RECT 17.110 2769.160 17.390 2769.440 ;
      LAYER met3 ;
        RECT -4.800 2769.450 2.400 2769.900 ;
        RECT 17.085 2769.450 17.415 2769.465 ;
        RECT -4.800 2769.150 17.415 2769.450 ;
        RECT -4.800 2768.700 2.400 2769.150 ;
        RECT 17.085 2769.135 17.415 2769.150 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 2505.020 15.570 2505.080 ;
        RECT 608.190 2505.020 608.510 2505.080 ;
        RECT 15.250 2504.880 608.510 2505.020 ;
        RECT 15.250 2504.820 15.570 2504.880 ;
        RECT 608.190 2504.820 608.510 2504.880 ;
      LAYER via ;
        RECT 15.280 2504.820 15.540 2505.080 ;
        RECT 608.220 2504.820 608.480 2505.080 ;
      LAYER met2 ;
        RECT 15.270 2508.675 15.550 2509.045 ;
        RECT 15.340 2505.110 15.480 2508.675 ;
        RECT 15.280 2504.790 15.540 2505.110 ;
        RECT 608.220 2504.790 608.480 2505.110 ;
        RECT 608.280 799.410 608.420 2504.790 ;
        RECT 609.390 799.410 609.670 800.000 ;
        RECT 608.280 799.270 609.670 799.410 ;
        RECT 609.390 796.000 609.670 799.270 ;
      LAYER via2 ;
        RECT 15.270 2508.720 15.550 2509.000 ;
      LAYER met3 ;
        RECT -4.800 2509.010 2.400 2509.460 ;
        RECT 15.245 2509.010 15.575 2509.025 ;
        RECT -4.800 2508.710 15.575 2509.010 ;
        RECT -4.800 2508.260 2.400 2508.710 ;
        RECT 15.245 2508.695 15.575 2508.710 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2242.880 16.030 2242.940 ;
        RECT 615.090 2242.880 615.410 2242.940 ;
        RECT 15.710 2242.740 615.410 2242.880 ;
        RECT 15.710 2242.680 16.030 2242.740 ;
        RECT 615.090 2242.680 615.410 2242.740 ;
      LAYER via ;
        RECT 15.740 2242.680 16.000 2242.940 ;
        RECT 615.120 2242.680 615.380 2242.940 ;
      LAYER met2 ;
        RECT 15.730 2247.555 16.010 2247.925 ;
        RECT 15.800 2242.970 15.940 2247.555 ;
        RECT 15.740 2242.650 16.000 2242.970 ;
        RECT 615.120 2242.650 615.380 2242.970 ;
        RECT 615.180 799.410 615.320 2242.650 ;
        RECT 616.290 799.410 616.570 800.000 ;
        RECT 615.180 799.270 616.570 799.410 ;
        RECT 616.290 796.000 616.570 799.270 ;
      LAYER via2 ;
        RECT 15.730 2247.600 16.010 2247.880 ;
      LAYER met3 ;
        RECT -4.800 2247.890 2.400 2248.340 ;
        RECT 15.705 2247.890 16.035 2247.905 ;
        RECT -4.800 2247.590 16.035 2247.890 ;
        RECT -4.800 2247.140 2.400 2247.590 ;
        RECT 15.705 2247.575 16.035 2247.590 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 1987.540 17.410 1987.600 ;
        RECT 621.990 1987.540 622.310 1987.600 ;
        RECT 17.090 1987.400 622.310 1987.540 ;
        RECT 17.090 1987.340 17.410 1987.400 ;
        RECT 621.990 1987.340 622.310 1987.400 ;
      LAYER via ;
        RECT 17.120 1987.340 17.380 1987.600 ;
        RECT 622.020 1987.340 622.280 1987.600 ;
      LAYER met2 ;
        RECT 17.120 1987.485 17.380 1987.630 ;
        RECT 17.110 1987.115 17.390 1987.485 ;
        RECT 622.020 1987.310 622.280 1987.630 ;
        RECT 622.080 799.410 622.220 1987.310 ;
        RECT 623.190 799.410 623.470 800.000 ;
        RECT 622.080 799.270 623.470 799.410 ;
        RECT 623.190 796.000 623.470 799.270 ;
      LAYER via2 ;
        RECT 17.110 1987.160 17.390 1987.440 ;
      LAYER met3 ;
        RECT -4.800 1987.450 2.400 1987.900 ;
        RECT 17.085 1987.450 17.415 1987.465 ;
        RECT -4.800 1987.150 17.415 1987.450 ;
        RECT -4.800 1986.700 2.400 1987.150 ;
        RECT 17.085 1987.135 17.415 1987.150 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 438.450 810.120 438.770 810.180 ;
        RECT 544.250 810.120 544.570 810.180 ;
        RECT 438.450 809.980 544.570 810.120 ;
        RECT 438.450 809.920 438.770 809.980 ;
        RECT 544.250 809.920 544.570 809.980 ;
        RECT 617.850 797.540 618.170 797.600 ;
        RECT 579.530 797.400 618.170 797.540 ;
        RECT 544.250 796.860 544.570 796.920 ;
        RECT 579.530 796.860 579.670 797.400 ;
        RECT 617.850 797.340 618.170 797.400 ;
        RECT 544.250 796.720 579.670 796.860 ;
        RECT 617.850 796.860 618.170 796.920 ;
        RECT 2903.590 796.860 2903.910 796.920 ;
        RECT 617.850 796.720 2903.910 796.860 ;
        RECT 544.250 796.660 544.570 796.720 ;
        RECT 617.850 796.660 618.170 796.720 ;
        RECT 2903.590 796.660 2903.910 796.720 ;
      LAYER via ;
        RECT 438.480 809.920 438.740 810.180 ;
        RECT 544.280 809.920 544.540 810.180 ;
        RECT 544.280 796.660 544.540 796.920 ;
        RECT 617.880 797.340 618.140 797.600 ;
        RECT 617.880 796.660 618.140 796.920 ;
        RECT 2903.620 796.660 2903.880 796.920 ;
      LAYER met2 ;
        RECT 438.480 809.890 438.740 810.210 ;
        RECT 544.280 809.890 544.540 810.210 ;
        RECT 436.890 799.410 437.170 800.000 ;
        RECT 438.540 799.410 438.680 809.890 ;
        RECT 436.890 799.270 438.680 799.410 ;
        RECT 436.890 796.000 437.170 799.270 ;
        RECT 544.340 796.950 544.480 809.890 ;
        RECT 617.880 797.310 618.140 797.630 ;
        RECT 617.940 796.950 618.080 797.310 ;
        RECT 544.280 796.630 544.540 796.950 ;
        RECT 617.880 796.630 618.140 796.950 ;
        RECT 2903.620 796.630 2903.880 796.950 ;
        RECT 2903.680 564.245 2903.820 796.630 ;
        RECT 2903.610 563.875 2903.890 564.245 ;
      LAYER via2 ;
        RECT 2903.610 563.920 2903.890 564.200 ;
      LAYER met3 ;
        RECT 2903.585 564.210 2903.915 564.225 ;
        RECT 2917.600 564.210 2924.800 564.660 ;
        RECT 2903.585 563.910 2924.800 564.210 ;
        RECT 2903.585 563.895 2903.915 563.910 ;
        RECT 2917.600 563.460 2924.800 563.910 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1725.400 16.950 1725.460 ;
        RECT 628.890 1725.400 629.210 1725.460 ;
        RECT 16.630 1725.260 629.210 1725.400 ;
        RECT 16.630 1725.200 16.950 1725.260 ;
        RECT 628.890 1725.200 629.210 1725.260 ;
      LAYER via ;
        RECT 16.660 1725.200 16.920 1725.460 ;
        RECT 628.920 1725.200 629.180 1725.460 ;
      LAYER met2 ;
        RECT 16.650 1726.675 16.930 1727.045 ;
        RECT 16.720 1725.490 16.860 1726.675 ;
        RECT 16.660 1725.170 16.920 1725.490 ;
        RECT 628.920 1725.170 629.180 1725.490 ;
        RECT 628.980 799.410 629.120 1725.170 ;
        RECT 630.090 799.410 630.370 800.000 ;
        RECT 628.980 799.270 630.370 799.410 ;
        RECT 630.090 796.000 630.370 799.270 ;
      LAYER via2 ;
        RECT 16.650 1726.720 16.930 1727.000 ;
      LAYER met3 ;
        RECT -4.800 1727.010 2.400 1727.460 ;
        RECT 16.625 1727.010 16.955 1727.025 ;
        RECT -4.800 1726.710 16.955 1727.010 ;
        RECT -4.800 1726.260 2.400 1726.710 ;
        RECT 16.625 1726.695 16.955 1726.710 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 1462.920 17.410 1462.980 ;
        RECT 635.790 1462.920 636.110 1462.980 ;
        RECT 17.090 1462.780 636.110 1462.920 ;
        RECT 17.090 1462.720 17.410 1462.780 ;
        RECT 635.790 1462.720 636.110 1462.780 ;
      LAYER via ;
        RECT 17.120 1462.720 17.380 1462.980 ;
        RECT 635.820 1462.720 636.080 1462.980 ;
      LAYER met2 ;
        RECT 17.110 1465.555 17.390 1465.925 ;
        RECT 17.180 1463.010 17.320 1465.555 ;
        RECT 17.120 1462.690 17.380 1463.010 ;
        RECT 635.820 1462.690 636.080 1463.010 ;
        RECT 635.880 799.410 636.020 1462.690 ;
        RECT 636.990 799.410 637.270 800.000 ;
        RECT 635.880 799.270 637.270 799.410 ;
        RECT 636.990 796.000 637.270 799.270 ;
      LAYER via2 ;
        RECT 17.110 1465.600 17.390 1465.880 ;
      LAYER met3 ;
        RECT -4.800 1465.890 2.400 1466.340 ;
        RECT 17.085 1465.890 17.415 1465.905 ;
        RECT -4.800 1465.590 17.415 1465.890 ;
        RECT -4.800 1465.140 2.400 1465.590 ;
        RECT 17.085 1465.575 17.415 1465.590 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 1200.780 17.410 1200.840 ;
        RECT 642.690 1200.780 643.010 1200.840 ;
        RECT 17.090 1200.640 643.010 1200.780 ;
        RECT 17.090 1200.580 17.410 1200.640 ;
        RECT 642.690 1200.580 643.010 1200.640 ;
      LAYER via ;
        RECT 17.120 1200.580 17.380 1200.840 ;
        RECT 642.720 1200.580 642.980 1200.840 ;
      LAYER met2 ;
        RECT 17.110 1205.115 17.390 1205.485 ;
        RECT 17.180 1200.870 17.320 1205.115 ;
        RECT 17.120 1200.550 17.380 1200.870 ;
        RECT 642.720 1200.550 642.980 1200.870 ;
        RECT 642.780 799.410 642.920 1200.550 ;
        RECT 643.890 799.410 644.170 800.000 ;
        RECT 642.780 799.270 644.170 799.410 ;
        RECT 643.890 796.000 644.170 799.270 ;
      LAYER via2 ;
        RECT 17.110 1205.160 17.390 1205.440 ;
      LAYER met3 ;
        RECT -4.800 1205.450 2.400 1205.900 ;
        RECT 17.085 1205.450 17.415 1205.465 ;
        RECT -4.800 1205.150 17.415 1205.450 ;
        RECT -4.800 1204.700 2.400 1205.150 ;
        RECT 17.085 1205.135 17.415 1205.150 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 938.640 17.410 938.700 ;
        RECT 649.590 938.640 649.910 938.700 ;
        RECT 17.090 938.500 649.910 938.640 ;
        RECT 17.090 938.440 17.410 938.500 ;
        RECT 649.590 938.440 649.910 938.500 ;
      LAYER via ;
        RECT 17.120 938.440 17.380 938.700 ;
        RECT 649.620 938.440 649.880 938.700 ;
      LAYER met2 ;
        RECT 17.110 943.995 17.390 944.365 ;
        RECT 17.180 938.730 17.320 943.995 ;
        RECT 17.120 938.410 17.380 938.730 ;
        RECT 649.620 938.410 649.880 938.730 ;
        RECT 649.680 799.410 649.820 938.410 ;
        RECT 650.790 799.410 651.070 800.000 ;
        RECT 649.680 799.270 651.070 799.410 ;
        RECT 650.790 796.000 651.070 799.270 ;
      LAYER via2 ;
        RECT 17.110 944.040 17.390 944.320 ;
      LAYER met3 ;
        RECT -4.800 944.330 2.400 944.780 ;
        RECT 17.085 944.330 17.415 944.345 ;
        RECT -4.800 944.030 17.415 944.330 ;
        RECT -4.800 943.580 2.400 944.030 ;
        RECT 17.085 944.015 17.415 944.030 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 37.790 808.420 38.110 808.480 ;
        RECT 656.030 808.420 656.350 808.480 ;
        RECT 37.790 808.280 656.350 808.420 ;
        RECT 37.790 808.220 38.110 808.280 ;
        RECT 656.030 808.220 656.350 808.280 ;
        RECT 14.330 688.400 14.650 688.460 ;
        RECT 37.790 688.400 38.110 688.460 ;
        RECT 14.330 688.260 38.110 688.400 ;
        RECT 14.330 688.200 14.650 688.260 ;
        RECT 37.790 688.200 38.110 688.260 ;
      LAYER via ;
        RECT 37.820 808.220 38.080 808.480 ;
        RECT 656.060 808.220 656.320 808.480 ;
        RECT 14.360 688.200 14.620 688.460 ;
        RECT 37.820 688.200 38.080 688.460 ;
      LAYER met2 ;
        RECT 37.820 808.190 38.080 808.510 ;
        RECT 656.060 808.190 656.320 808.510 ;
        RECT 37.880 688.490 38.020 808.190 ;
        RECT 656.120 799.410 656.260 808.190 ;
        RECT 657.690 799.410 657.970 800.000 ;
        RECT 656.120 799.270 657.970 799.410 ;
        RECT 657.690 796.000 657.970 799.270 ;
        RECT 14.360 688.170 14.620 688.490 ;
        RECT 37.820 688.170 38.080 688.490 ;
        RECT 14.420 683.925 14.560 688.170 ;
        RECT 14.350 683.555 14.630 683.925 ;
      LAYER via2 ;
        RECT 14.350 683.600 14.630 683.880 ;
      LAYER met3 ;
        RECT -4.800 683.890 2.400 684.340 ;
        RECT 14.325 683.890 14.655 683.905 ;
        RECT -4.800 683.590 14.655 683.890 ;
        RECT -4.800 683.140 2.400 683.590 ;
        RECT 14.325 683.575 14.655 683.590 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 663.390 797.200 663.710 797.260 ;
        RECT 420.830 797.060 469.270 797.200 ;
        RECT 417.290 793.800 417.610 793.860 ;
        RECT 420.830 793.800 420.970 797.060 ;
        RECT 469.130 795.500 469.270 797.060 ;
        RECT 604.140 797.060 663.710 797.200 ;
        RECT 469.130 795.360 476.170 795.500 ;
        RECT 476.030 795.160 476.170 795.360 ;
        RECT 476.030 795.020 483.070 795.160 ;
        RECT 482.930 794.480 483.070 795.020 ;
        RECT 604.140 794.480 604.280 797.060 ;
        RECT 663.390 797.000 663.710 797.060 ;
        RECT 482.930 794.340 604.280 794.480 ;
        RECT 417.290 793.660 420.970 793.800 ;
        RECT 417.290 793.600 417.610 793.660 ;
        RECT 15.710 427.620 16.030 427.680 ;
        RECT 417.290 427.620 417.610 427.680 ;
        RECT 15.710 427.480 417.610 427.620 ;
        RECT 15.710 427.420 16.030 427.480 ;
        RECT 417.290 427.420 417.610 427.480 ;
      LAYER via ;
        RECT 417.320 793.600 417.580 793.860 ;
        RECT 663.420 797.000 663.680 797.260 ;
        RECT 15.740 427.420 16.000 427.680 ;
        RECT 417.320 427.420 417.580 427.680 ;
      LAYER met2 ;
        RECT 664.590 797.370 664.870 800.000 ;
        RECT 663.480 797.290 664.870 797.370 ;
        RECT 663.420 797.230 664.870 797.290 ;
        RECT 663.420 796.970 663.680 797.230 ;
        RECT 664.590 796.000 664.870 797.230 ;
        RECT 417.320 793.570 417.580 793.890 ;
        RECT 417.380 427.710 417.520 793.570 ;
        RECT 15.740 427.390 16.000 427.710 ;
        RECT 417.320 427.390 417.580 427.710 ;
        RECT 15.800 423.485 15.940 427.390 ;
        RECT 15.730 423.115 16.010 423.485 ;
      LAYER via2 ;
        RECT 15.730 423.160 16.010 423.440 ;
      LAYER met3 ;
        RECT -4.800 423.450 2.400 423.900 ;
        RECT 15.705 423.450 16.035 423.465 ;
        RECT -4.800 423.150 16.035 423.450 ;
        RECT -4.800 422.700 2.400 423.150 ;
        RECT 15.705 423.135 16.035 423.150 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 802.300 17.870 802.360 ;
        RECT 669.830 802.300 670.150 802.360 ;
        RECT 17.550 802.160 670.150 802.300 ;
        RECT 17.550 802.100 17.870 802.160 ;
        RECT 669.830 802.100 670.150 802.160 ;
      LAYER via ;
        RECT 17.580 802.100 17.840 802.360 ;
        RECT 669.860 802.100 670.120 802.360 ;
      LAYER met2 ;
        RECT 17.580 802.070 17.840 802.390 ;
        RECT 669.860 802.070 670.120 802.390 ;
        RECT 17.640 227.645 17.780 802.070 ;
        RECT 669.920 799.410 670.060 802.070 ;
        RECT 671.490 799.410 671.770 800.000 ;
        RECT 669.920 799.270 671.770 799.410 ;
        RECT 671.490 796.000 671.770 799.270 ;
        RECT 17.570 227.275 17.850 227.645 ;
      LAYER via2 ;
        RECT 17.570 227.320 17.850 227.600 ;
      LAYER met3 ;
        RECT -4.800 227.610 2.400 228.060 ;
        RECT 17.545 227.610 17.875 227.625 ;
        RECT -4.800 227.310 17.875 227.610 ;
        RECT -4.800 226.860 2.400 227.310 ;
        RECT 17.545 227.295 17.875 227.310 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 34.240 17.410 34.300 ;
        RECT 681.330 34.240 681.650 34.300 ;
        RECT 17.090 34.100 681.650 34.240 ;
        RECT 17.090 34.040 17.410 34.100 ;
        RECT 681.330 34.040 681.650 34.100 ;
      LAYER via ;
        RECT 17.120 34.040 17.380 34.300 ;
        RECT 681.360 34.040 681.620 34.300 ;
      LAYER met2 ;
        RECT 678.390 796.690 678.670 800.000 ;
        RECT 679.510 796.690 679.790 796.805 ;
        RECT 678.390 796.550 679.790 796.690 ;
        RECT 678.390 796.000 678.670 796.550 ;
        RECT 679.510 796.435 679.790 796.550 ;
        RECT 681.350 795.755 681.630 796.125 ;
        RECT 681.420 34.330 681.560 795.755 ;
        RECT 17.120 34.010 17.380 34.330 ;
        RECT 681.360 34.010 681.620 34.330 ;
        RECT 17.180 32.485 17.320 34.010 ;
        RECT 17.110 32.115 17.390 32.485 ;
      LAYER via2 ;
        RECT 679.510 796.480 679.790 796.760 ;
        RECT 681.350 795.800 681.630 796.080 ;
        RECT 17.110 32.160 17.390 32.440 ;
      LAYER met3 ;
        RECT 679.485 796.770 679.815 796.785 ;
        RECT 679.485 796.470 681.410 796.770 ;
        RECT 679.485 796.455 679.815 796.470 ;
        RECT 681.110 796.105 681.410 796.470 ;
        RECT 681.110 795.790 681.655 796.105 ;
        RECT 681.325 795.775 681.655 795.790 ;
        RECT -4.800 32.450 2.400 32.900 ;
        RECT 17.085 32.450 17.415 32.465 ;
        RECT -4.800 32.150 17.415 32.450 ;
        RECT -4.800 31.700 2.400 32.150 ;
        RECT 17.085 32.135 17.415 32.150 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 445.350 807.400 445.670 807.460 ;
        RECT 2904.510 807.400 2904.830 807.460 ;
        RECT 445.350 807.260 2904.830 807.400 ;
        RECT 445.350 807.200 445.670 807.260 ;
        RECT 2904.510 807.200 2904.830 807.260 ;
      LAYER via ;
        RECT 445.380 807.200 445.640 807.460 ;
        RECT 2904.540 807.200 2904.800 807.460 ;
      LAYER met2 ;
        RECT 445.380 807.170 445.640 807.490 ;
        RECT 2904.540 807.170 2904.800 807.490 ;
        RECT 443.790 799.410 444.070 800.000 ;
        RECT 445.440 799.410 445.580 807.170 ;
        RECT 443.790 799.270 445.580 799.410 ;
        RECT 443.790 796.000 444.070 799.270 ;
        RECT 2904.600 763.485 2904.740 807.170 ;
        RECT 2904.530 763.115 2904.810 763.485 ;
      LAYER via2 ;
        RECT 2904.530 763.160 2904.810 763.440 ;
      LAYER met3 ;
        RECT 2904.505 763.450 2904.835 763.465 ;
        RECT 2917.600 763.450 2924.800 763.900 ;
        RECT 2904.505 763.150 2924.800 763.450 ;
        RECT 2904.505 763.135 2904.835 763.150 ;
        RECT 2917.600 762.700 2924.800 763.150 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 449.030 959.380 449.350 959.440 ;
        RECT 2900.830 959.380 2901.150 959.440 ;
        RECT 449.030 959.240 2901.150 959.380 ;
        RECT 449.030 959.180 449.350 959.240 ;
        RECT 2900.830 959.180 2901.150 959.240 ;
      LAYER via ;
        RECT 449.060 959.180 449.320 959.440 ;
        RECT 2900.860 959.180 2901.120 959.440 ;
      LAYER met2 ;
        RECT 2900.850 962.355 2901.130 962.725 ;
        RECT 2900.920 959.470 2901.060 962.355 ;
        RECT 449.060 959.150 449.320 959.470 ;
        RECT 2900.860 959.150 2901.120 959.470 ;
        RECT 449.120 799.410 449.260 959.150 ;
        RECT 450.690 799.410 450.970 800.000 ;
        RECT 449.120 799.270 450.970 799.410 ;
        RECT 450.690 796.000 450.970 799.270 ;
      LAYER via2 ;
        RECT 2900.850 962.400 2901.130 962.680 ;
      LAYER met3 ;
        RECT 2900.825 962.690 2901.155 962.705 ;
        RECT 2917.600 962.690 2924.800 963.140 ;
        RECT 2900.825 962.390 2924.800 962.690 ;
        RECT 2900.825 962.375 2901.155 962.390 ;
        RECT 2917.600 961.940 2924.800 962.390 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.930 1159.300 456.250 1159.360 ;
        RECT 2900.830 1159.300 2901.150 1159.360 ;
        RECT 455.930 1159.160 2901.150 1159.300 ;
        RECT 455.930 1159.100 456.250 1159.160 ;
        RECT 2900.830 1159.100 2901.150 1159.160 ;
      LAYER via ;
        RECT 455.960 1159.100 456.220 1159.360 ;
        RECT 2900.860 1159.100 2901.120 1159.360 ;
      LAYER met2 ;
        RECT 2900.850 1161.595 2901.130 1161.965 ;
        RECT 2900.920 1159.390 2901.060 1161.595 ;
        RECT 455.960 1159.070 456.220 1159.390 ;
        RECT 2900.860 1159.070 2901.120 1159.390 ;
        RECT 456.020 799.410 456.160 1159.070 ;
        RECT 457.590 799.410 457.870 800.000 ;
        RECT 456.020 799.270 457.870 799.410 ;
        RECT 457.590 796.000 457.870 799.270 ;
      LAYER via2 ;
        RECT 2900.850 1161.640 2901.130 1161.920 ;
      LAYER met3 ;
        RECT 2900.825 1161.930 2901.155 1161.945 ;
        RECT 2917.600 1161.930 2924.800 1162.380 ;
        RECT 2900.825 1161.630 2924.800 1161.930 ;
        RECT 2900.825 1161.615 2901.155 1161.630 ;
        RECT 2917.600 1161.180 2924.800 1161.630 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.830 1359.560 463.150 1359.620 ;
        RECT 2898.990 1359.560 2899.310 1359.620 ;
        RECT 462.830 1359.420 2899.310 1359.560 ;
        RECT 462.830 1359.360 463.150 1359.420 ;
        RECT 2898.990 1359.360 2899.310 1359.420 ;
      LAYER via ;
        RECT 462.860 1359.360 463.120 1359.620 ;
        RECT 2899.020 1359.360 2899.280 1359.620 ;
      LAYER met2 ;
        RECT 2899.010 1360.835 2899.290 1361.205 ;
        RECT 2899.080 1359.650 2899.220 1360.835 ;
        RECT 462.860 1359.330 463.120 1359.650 ;
        RECT 2899.020 1359.330 2899.280 1359.650 ;
        RECT 462.920 799.410 463.060 1359.330 ;
        RECT 464.490 799.410 464.770 800.000 ;
        RECT 462.920 799.270 464.770 799.410 ;
        RECT 464.490 796.000 464.770 799.270 ;
      LAYER via2 ;
        RECT 2899.010 1360.880 2899.290 1361.160 ;
      LAYER met3 ;
        RECT 2898.985 1361.170 2899.315 1361.185 ;
        RECT 2917.600 1361.170 2924.800 1361.620 ;
        RECT 2898.985 1360.870 2924.800 1361.170 ;
        RECT 2898.985 1360.855 2899.315 1360.870 ;
        RECT 2917.600 1360.420 2924.800 1360.870 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.730 1621.700 470.050 1621.760 ;
        RECT 2900.830 1621.700 2901.150 1621.760 ;
        RECT 469.730 1621.560 2901.150 1621.700 ;
        RECT 469.730 1621.500 470.050 1621.560 ;
        RECT 2900.830 1621.500 2901.150 1621.560 ;
      LAYER via ;
        RECT 469.760 1621.500 470.020 1621.760 ;
        RECT 2900.860 1621.500 2901.120 1621.760 ;
      LAYER met2 ;
        RECT 2900.850 1626.035 2901.130 1626.405 ;
        RECT 2900.920 1621.790 2901.060 1626.035 ;
        RECT 469.760 1621.470 470.020 1621.790 ;
        RECT 2900.860 1621.470 2901.120 1621.790 ;
        RECT 469.820 799.410 469.960 1621.470 ;
        RECT 471.390 799.410 471.670 800.000 ;
        RECT 469.820 799.270 471.670 799.410 ;
        RECT 471.390 796.000 471.670 799.270 ;
      LAYER via2 ;
        RECT 2900.850 1626.080 2901.130 1626.360 ;
      LAYER met3 ;
        RECT 2900.825 1626.370 2901.155 1626.385 ;
        RECT 2917.600 1626.370 2924.800 1626.820 ;
        RECT 2900.825 1626.070 2924.800 1626.370 ;
        RECT 2900.825 1626.055 2901.155 1626.070 ;
        RECT 2917.600 1625.620 2924.800 1626.070 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.630 1890.980 476.950 1891.040 ;
        RECT 2900.830 1890.980 2901.150 1891.040 ;
        RECT 476.630 1890.840 2901.150 1890.980 ;
        RECT 476.630 1890.780 476.950 1890.840 ;
        RECT 2900.830 1890.780 2901.150 1890.840 ;
      LAYER via ;
        RECT 476.660 1890.780 476.920 1891.040 ;
        RECT 2900.860 1890.780 2901.120 1891.040 ;
      LAYER met2 ;
        RECT 2900.850 1891.915 2901.130 1892.285 ;
        RECT 2900.920 1891.070 2901.060 1891.915 ;
        RECT 476.660 1890.750 476.920 1891.070 ;
        RECT 2900.860 1890.750 2901.120 1891.070 ;
        RECT 476.720 799.410 476.860 1890.750 ;
        RECT 478.290 799.410 478.570 800.000 ;
        RECT 476.720 799.270 478.570 799.410 ;
        RECT 478.290 796.000 478.570 799.270 ;
      LAYER via2 ;
        RECT 2900.850 1891.960 2901.130 1892.240 ;
      LAYER met3 ;
        RECT 2900.825 1892.250 2901.155 1892.265 ;
        RECT 2917.600 1892.250 2924.800 1892.700 ;
        RECT 2900.825 1891.950 2924.800 1892.250 ;
        RECT 2900.825 1891.935 2901.155 1891.950 ;
        RECT 2917.600 1891.500 2924.800 1891.950 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.530 2153.120 483.850 2153.180 ;
        RECT 2900.830 2153.120 2901.150 2153.180 ;
        RECT 483.530 2152.980 2901.150 2153.120 ;
        RECT 483.530 2152.920 483.850 2152.980 ;
        RECT 2900.830 2152.920 2901.150 2152.980 ;
      LAYER via ;
        RECT 483.560 2152.920 483.820 2153.180 ;
        RECT 2900.860 2152.920 2901.120 2153.180 ;
      LAYER met2 ;
        RECT 2900.850 2157.795 2901.130 2158.165 ;
        RECT 2900.920 2153.210 2901.060 2157.795 ;
        RECT 483.560 2152.890 483.820 2153.210 ;
        RECT 2900.860 2152.890 2901.120 2153.210 ;
        RECT 483.620 799.410 483.760 2152.890 ;
        RECT 485.190 799.410 485.470 800.000 ;
        RECT 483.620 799.270 485.470 799.410 ;
        RECT 485.190 796.000 485.470 799.270 ;
      LAYER via2 ;
        RECT 2900.850 2157.840 2901.130 2158.120 ;
      LAYER met3 ;
        RECT 2900.825 2158.130 2901.155 2158.145 ;
        RECT 2917.600 2158.130 2924.800 2158.580 ;
        RECT 2900.825 2157.830 2924.800 2158.130 ;
        RECT 2900.825 2157.815 2901.155 2157.830 ;
        RECT 2917.600 2157.380 2924.800 2157.830 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 426.950 807.740 427.270 807.800 ;
        RECT 1259.090 807.740 1259.410 807.800 ;
        RECT 426.950 807.600 1259.410 807.740 ;
        RECT 426.950 807.540 427.270 807.600 ;
        RECT 1259.090 807.540 1259.410 807.600 ;
        RECT 1259.090 107.680 1259.410 107.740 ;
        RECT 2900.830 107.680 2901.150 107.740 ;
        RECT 1259.090 107.540 2901.150 107.680 ;
        RECT 1259.090 107.480 1259.410 107.540 ;
        RECT 2900.830 107.480 2901.150 107.540 ;
      LAYER via ;
        RECT 426.980 807.540 427.240 807.800 ;
        RECT 1259.120 807.540 1259.380 807.800 ;
        RECT 1259.120 107.480 1259.380 107.740 ;
        RECT 2900.860 107.480 2901.120 107.740 ;
      LAYER met2 ;
        RECT 426.980 807.510 427.240 807.830 ;
        RECT 1259.120 807.510 1259.380 807.830 ;
        RECT 425.390 799.410 425.670 800.000 ;
        RECT 427.040 799.410 427.180 807.510 ;
        RECT 425.390 799.270 427.180 799.410 ;
        RECT 425.390 796.000 425.670 799.270 ;
        RECT 1259.180 107.770 1259.320 807.510 ;
        RECT 1259.120 107.450 1259.380 107.770 ;
        RECT 2900.860 107.450 2901.120 107.770 ;
        RECT 2900.920 99.125 2901.060 107.450 ;
        RECT 2900.850 98.755 2901.130 99.125 ;
      LAYER via2 ;
        RECT 2900.850 98.800 2901.130 99.080 ;
      LAYER met3 ;
        RECT 2900.825 99.090 2901.155 99.105 ;
        RECT 2917.600 99.090 2924.800 99.540 ;
        RECT 2900.825 98.790 2924.800 99.090 ;
        RECT 2900.825 98.775 2901.155 98.790 ;
        RECT 2917.600 98.340 2924.800 98.790 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.890 2353.040 491.210 2353.100 ;
        RECT 2899.910 2353.040 2900.230 2353.100 ;
        RECT 490.890 2352.900 2900.230 2353.040 ;
        RECT 490.890 2352.840 491.210 2352.900 ;
        RECT 2899.910 2352.840 2900.230 2352.900 ;
      LAYER via ;
        RECT 490.920 2352.840 491.180 2353.100 ;
        RECT 2899.940 2352.840 2900.200 2353.100 ;
      LAYER met2 ;
        RECT 2899.930 2357.035 2900.210 2357.405 ;
        RECT 2900.000 2353.130 2900.140 2357.035 ;
        RECT 490.920 2352.810 491.180 2353.130 ;
        RECT 2899.940 2352.810 2900.200 2353.130 ;
        RECT 490.980 855.670 491.120 2352.810 ;
        RECT 490.980 855.530 492.960 855.670 ;
        RECT 492.820 799.410 492.960 855.530 ;
        RECT 494.390 799.410 494.670 800.000 ;
        RECT 492.820 799.270 494.670 799.410 ;
        RECT 494.390 796.000 494.670 799.270 ;
      LAYER via2 ;
        RECT 2899.930 2357.080 2900.210 2357.360 ;
      LAYER met3 ;
        RECT 2899.905 2357.370 2900.235 2357.385 ;
        RECT 2917.600 2357.370 2924.800 2357.820 ;
        RECT 2899.905 2357.070 2924.800 2357.370 ;
        RECT 2899.905 2357.055 2900.235 2357.070 ;
        RECT 2917.600 2356.620 2924.800 2357.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.790 2622.320 498.110 2622.380 ;
        RECT 2900.830 2622.320 2901.150 2622.380 ;
        RECT 497.790 2622.180 2901.150 2622.320 ;
        RECT 497.790 2622.120 498.110 2622.180 ;
        RECT 2900.830 2622.120 2901.150 2622.180 ;
      LAYER via ;
        RECT 497.820 2622.120 498.080 2622.380 ;
        RECT 2900.860 2622.120 2901.120 2622.380 ;
      LAYER met2 ;
        RECT 497.820 2622.090 498.080 2622.410 ;
        RECT 2900.850 2622.235 2901.130 2622.605 ;
        RECT 2900.860 2622.090 2901.120 2622.235 ;
        RECT 497.880 855.670 498.020 2622.090 ;
        RECT 497.880 855.530 499.860 855.670 ;
        RECT 499.720 799.410 499.860 855.530 ;
        RECT 501.290 799.410 501.570 800.000 ;
        RECT 499.720 799.270 501.570 799.410 ;
        RECT 501.290 796.000 501.570 799.270 ;
      LAYER via2 ;
        RECT 2900.850 2622.280 2901.130 2622.560 ;
      LAYER met3 ;
        RECT 2900.825 2622.570 2901.155 2622.585 ;
        RECT 2917.600 2622.570 2924.800 2623.020 ;
        RECT 2900.825 2622.270 2924.800 2622.570 ;
        RECT 2900.825 2622.255 2901.155 2622.270 ;
        RECT 2917.600 2621.820 2924.800 2622.270 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.690 2884.460 505.010 2884.520 ;
        RECT 2900.830 2884.460 2901.150 2884.520 ;
        RECT 504.690 2884.320 2901.150 2884.460 ;
        RECT 504.690 2884.260 505.010 2884.320 ;
        RECT 2900.830 2884.260 2901.150 2884.320 ;
      LAYER via ;
        RECT 504.720 2884.260 504.980 2884.520 ;
        RECT 2900.860 2884.260 2901.120 2884.520 ;
      LAYER met2 ;
        RECT 2900.850 2888.115 2901.130 2888.485 ;
        RECT 2900.920 2884.550 2901.060 2888.115 ;
        RECT 504.720 2884.230 504.980 2884.550 ;
        RECT 2900.860 2884.230 2901.120 2884.550 ;
        RECT 504.780 855.670 504.920 2884.230 ;
        RECT 504.780 855.530 506.760 855.670 ;
        RECT 506.620 799.410 506.760 855.530 ;
        RECT 508.190 799.410 508.470 800.000 ;
        RECT 506.620 799.270 508.470 799.410 ;
        RECT 508.190 796.000 508.470 799.270 ;
      LAYER via2 ;
        RECT 2900.850 2888.160 2901.130 2888.440 ;
      LAYER met3 ;
        RECT 2900.825 2888.450 2901.155 2888.465 ;
        RECT 2917.600 2888.450 2924.800 2888.900 ;
        RECT 2900.825 2888.150 2924.800 2888.450 ;
        RECT 2900.825 2888.135 2901.155 2888.150 ;
        RECT 2917.600 2887.700 2924.800 2888.150 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.590 3153.400 511.910 3153.460 ;
        RECT 2900.830 3153.400 2901.150 3153.460 ;
        RECT 511.590 3153.260 2901.150 3153.400 ;
        RECT 511.590 3153.200 511.910 3153.260 ;
        RECT 2900.830 3153.200 2901.150 3153.260 ;
      LAYER via ;
        RECT 511.620 3153.200 511.880 3153.460 ;
        RECT 2900.860 3153.200 2901.120 3153.460 ;
      LAYER met2 ;
        RECT 2900.850 3153.995 2901.130 3154.365 ;
        RECT 2900.920 3153.490 2901.060 3153.995 ;
        RECT 511.620 3153.170 511.880 3153.490 ;
        RECT 2900.860 3153.170 2901.120 3153.490 ;
        RECT 511.680 855.670 511.820 3153.170 ;
        RECT 511.680 855.530 513.660 855.670 ;
        RECT 513.520 799.410 513.660 855.530 ;
        RECT 515.090 799.410 515.370 800.000 ;
        RECT 513.520 799.270 515.370 799.410 ;
        RECT 515.090 796.000 515.370 799.270 ;
      LAYER via2 ;
        RECT 2900.850 3154.040 2901.130 3154.320 ;
      LAYER met3 ;
        RECT 2900.825 3154.330 2901.155 3154.345 ;
        RECT 2917.600 3154.330 2924.800 3154.780 ;
        RECT 2900.825 3154.030 2924.800 3154.330 ;
        RECT 2900.825 3154.015 2901.155 3154.030 ;
        RECT 2917.600 3153.580 2924.800 3154.030 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.490 3415.880 518.810 3415.940 ;
        RECT 2900.830 3415.880 2901.150 3415.940 ;
        RECT 518.490 3415.740 2901.150 3415.880 ;
        RECT 518.490 3415.680 518.810 3415.740 ;
        RECT 2900.830 3415.680 2901.150 3415.740 ;
      LAYER via ;
        RECT 518.520 3415.680 518.780 3415.940 ;
        RECT 2900.860 3415.680 2901.120 3415.940 ;
      LAYER met2 ;
        RECT 2900.850 3419.195 2901.130 3419.565 ;
        RECT 2900.920 3415.970 2901.060 3419.195 ;
        RECT 518.520 3415.650 518.780 3415.970 ;
        RECT 2900.860 3415.650 2901.120 3415.970 ;
        RECT 518.580 855.670 518.720 3415.650 ;
        RECT 518.580 855.530 520.560 855.670 ;
        RECT 520.420 799.410 520.560 855.530 ;
        RECT 521.990 799.410 522.270 800.000 ;
        RECT 520.420 799.270 522.270 799.410 ;
        RECT 521.990 796.000 522.270 799.270 ;
      LAYER via2 ;
        RECT 2900.850 3419.240 2901.130 3419.520 ;
      LAYER met3 ;
        RECT 2900.825 3419.530 2901.155 3419.545 ;
        RECT 2917.600 3419.530 2924.800 3419.980 ;
        RECT 2900.825 3419.230 2924.800 3419.530 ;
        RECT 2900.825 3419.215 2901.155 3419.230 ;
        RECT 2917.600 3418.780 2924.800 3419.230 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 534.590 3501.560 534.910 3501.620 ;
        RECT 2717.290 3501.560 2717.610 3501.620 ;
        RECT 534.590 3501.420 2717.610 3501.560 ;
        RECT 534.590 3501.360 534.910 3501.420 ;
        RECT 2717.290 3501.360 2717.610 3501.420 ;
        RECT 529.990 814.200 530.310 814.260 ;
        RECT 534.590 814.200 534.910 814.260 ;
        RECT 529.990 814.060 534.910 814.200 ;
        RECT 529.990 814.000 530.310 814.060 ;
        RECT 534.590 814.000 534.910 814.060 ;
      LAYER via ;
        RECT 534.620 3501.360 534.880 3501.620 ;
        RECT 2717.320 3501.360 2717.580 3501.620 ;
        RECT 530.020 814.000 530.280 814.260 ;
        RECT 534.620 814.000 534.880 814.260 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.650 2717.520 3517.600 ;
        RECT 534.620 3501.330 534.880 3501.650 ;
        RECT 2717.320 3501.330 2717.580 3501.650 ;
        RECT 534.680 814.290 534.820 3501.330 ;
        RECT 530.020 813.970 530.280 814.290 ;
        RECT 534.620 813.970 534.880 814.290 ;
        RECT 528.890 799.410 529.170 800.000 ;
        RECT 530.080 799.410 530.220 813.970 ;
        RECT 528.890 799.270 530.220 799.410 ;
        RECT 528.890 796.000 529.170 799.270 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.830 831.540 532.150 831.600 ;
        RECT 2387.470 831.540 2387.790 831.600 ;
        RECT 531.830 831.400 2387.790 831.540 ;
        RECT 531.830 831.340 532.150 831.400 ;
        RECT 2387.470 831.340 2387.790 831.400 ;
        RECT 531.830 803.660 532.150 803.720 ;
        RECT 534.130 803.660 534.450 803.720 ;
        RECT 531.830 803.520 534.450 803.660 ;
        RECT 531.830 803.460 532.150 803.520 ;
        RECT 534.130 803.460 534.450 803.520 ;
      LAYER via ;
        RECT 531.860 831.340 532.120 831.600 ;
        RECT 2387.500 831.340 2387.760 831.600 ;
        RECT 531.860 803.460 532.120 803.720 ;
        RECT 534.160 803.460 534.420 803.720 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3512.170 2392.760 3517.600 ;
        RECT 2387.560 3512.030 2392.760 3512.170 ;
        RECT 2387.560 831.630 2387.700 3512.030 ;
        RECT 531.860 831.310 532.120 831.630 ;
        RECT 2387.500 831.310 2387.760 831.630 ;
        RECT 531.920 803.750 532.060 831.310 ;
        RECT 531.860 803.430 532.120 803.750 ;
        RECT 534.160 803.430 534.420 803.750 ;
        RECT 534.220 799.410 534.360 803.430 ;
        RECT 535.790 799.410 536.070 800.000 ;
        RECT 534.220 799.270 536.070 799.410 ;
        RECT 535.790 796.000 536.070 799.270 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.730 3501.900 539.050 3501.960 ;
        RECT 2068.230 3501.900 2068.550 3501.960 ;
        RECT 538.730 3501.760 2068.550 3501.900 ;
        RECT 538.730 3501.700 539.050 3501.760 ;
        RECT 2068.230 3501.700 2068.550 3501.760 ;
      LAYER via ;
        RECT 538.760 3501.700 539.020 3501.960 ;
        RECT 2068.260 3501.700 2068.520 3501.960 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3501.990 2068.460 3517.600 ;
        RECT 538.760 3501.670 539.020 3501.990 ;
        RECT 2068.260 3501.670 2068.520 3501.990 ;
        RECT 538.820 855.670 538.960 3501.670 ;
        RECT 538.820 855.530 541.260 855.670 ;
        RECT 541.120 799.410 541.260 855.530 ;
        RECT 542.690 799.410 542.970 800.000 ;
        RECT 541.120 799.270 542.970 799.410 ;
        RECT 542.690 796.000 542.970 799.270 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 693.290 3502.240 693.610 3502.300 ;
        RECT 1743.930 3502.240 1744.250 3502.300 ;
        RECT 693.290 3502.100 1744.250 3502.240 ;
        RECT 693.290 3502.040 693.610 3502.100 ;
        RECT 1743.930 3502.040 1744.250 3502.100 ;
        RECT 551.150 810.800 551.470 810.860 ;
        RECT 693.290 810.800 693.610 810.860 ;
        RECT 551.150 810.660 693.610 810.800 ;
        RECT 551.150 810.600 551.470 810.660 ;
        RECT 693.290 810.600 693.610 810.660 ;
      LAYER via ;
        RECT 693.320 3502.040 693.580 3502.300 ;
        RECT 1743.960 3502.040 1744.220 3502.300 ;
        RECT 551.180 810.600 551.440 810.860 ;
        RECT 693.320 810.600 693.580 810.860 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3502.330 1744.160 3517.600 ;
        RECT 693.320 3502.010 693.580 3502.330 ;
        RECT 1743.960 3502.010 1744.220 3502.330 ;
        RECT 693.380 810.890 693.520 3502.010 ;
        RECT 551.180 810.570 551.440 810.890 ;
        RECT 693.320 810.570 693.580 810.890 ;
        RECT 549.590 799.410 549.870 800.000 ;
        RECT 551.240 799.410 551.380 810.570 ;
        RECT 549.590 799.270 551.380 799.410 ;
        RECT 549.590 796.000 549.870 799.270 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.530 3502.580 552.850 3502.640 ;
        RECT 1419.170 3502.580 1419.490 3502.640 ;
        RECT 552.530 3502.440 1419.490 3502.580 ;
        RECT 552.530 3502.380 552.850 3502.440 ;
        RECT 1419.170 3502.380 1419.490 3502.440 ;
      LAYER via ;
        RECT 552.560 3502.380 552.820 3502.640 ;
        RECT 1419.200 3502.380 1419.460 3502.640 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3502.670 1419.400 3517.600 ;
        RECT 552.560 3502.350 552.820 3502.670 ;
        RECT 1419.200 3502.350 1419.460 3502.670 ;
        RECT 552.620 855.670 552.760 3502.350 ;
        RECT 552.620 855.530 555.060 855.670 ;
        RECT 554.920 799.410 555.060 855.530 ;
        RECT 556.490 799.410 556.770 800.000 ;
        RECT 554.920 799.270 556.770 799.410 ;
        RECT 556.490 796.000 556.770 799.270 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.790 810.120 567.110 810.180 ;
        RECT 565.730 809.980 567.110 810.120 ;
        RECT 433.850 809.780 434.170 809.840 ;
        RECT 565.730 809.780 565.870 809.980 ;
        RECT 566.790 809.920 567.110 809.980 ;
        RECT 433.850 809.640 565.870 809.780 ;
        RECT 433.850 809.580 434.170 809.640 ;
        RECT 566.790 803.660 567.110 803.720 ;
        RECT 2902.670 803.660 2902.990 803.720 ;
        RECT 566.790 803.520 2902.990 803.660 ;
        RECT 566.790 803.460 567.110 803.520 ;
        RECT 2902.670 803.460 2902.990 803.520 ;
      LAYER via ;
        RECT 433.880 809.580 434.140 809.840 ;
        RECT 566.820 809.920 567.080 810.180 ;
        RECT 566.820 803.460 567.080 803.720 ;
        RECT 2902.700 803.460 2902.960 803.720 ;
      LAYER met2 ;
        RECT 566.820 809.890 567.080 810.210 ;
        RECT 433.880 809.550 434.140 809.870 ;
        RECT 432.290 799.410 432.570 800.000 ;
        RECT 433.940 799.410 434.080 809.550 ;
        RECT 566.880 803.750 567.020 809.890 ;
        RECT 566.820 803.430 567.080 803.750 ;
        RECT 2902.700 803.430 2902.960 803.750 ;
        RECT 432.290 799.270 434.080 799.410 ;
        RECT 432.290 796.000 432.570 799.270 ;
        RECT 2902.760 298.365 2902.900 803.430 ;
        RECT 2902.690 297.995 2902.970 298.365 ;
      LAYER via2 ;
        RECT 2902.690 298.040 2902.970 298.320 ;
      LAYER met3 ;
        RECT 2902.665 298.330 2902.995 298.345 ;
        RECT 2917.600 298.330 2924.800 298.780 ;
        RECT 2902.665 298.030 2924.800 298.330 ;
        RECT 2902.665 298.015 2902.995 298.030 ;
        RECT 2917.600 297.580 2924.800 298.030 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 561.730 832.220 562.050 832.280 ;
        RECT 1090.270 832.220 1090.590 832.280 ;
        RECT 561.730 832.080 1090.590 832.220 ;
        RECT 561.730 832.020 562.050 832.080 ;
        RECT 1090.270 832.020 1090.590 832.080 ;
      LAYER via ;
        RECT 561.760 832.020 562.020 832.280 ;
        RECT 1090.300 832.020 1090.560 832.280 ;
      LAYER met2 ;
        RECT 1090.360 3517.910 1094.180 3518.050 ;
        RECT 1090.360 832.310 1090.500 3517.910 ;
        RECT 1094.040 3517.370 1094.180 3517.910 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3517.370 1095.100 3517.600 ;
        RECT 1094.040 3517.230 1095.100 3517.370 ;
        RECT 561.760 831.990 562.020 832.310 ;
        RECT 1090.300 831.990 1090.560 832.310 ;
        RECT 561.820 799.410 561.960 831.990 ;
        RECT 563.390 799.410 563.670 800.000 ;
        RECT 561.820 799.270 563.670 799.410 ;
        RECT 563.390 796.000 563.670 799.270 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 700.190 3503.260 700.510 3503.320 ;
        RECT 770.570 3503.260 770.890 3503.320 ;
        RECT 700.190 3503.120 770.890 3503.260 ;
        RECT 700.190 3503.060 700.510 3503.120 ;
        RECT 770.570 3503.060 770.890 3503.120 ;
        RECT 571.850 811.140 572.170 811.200 ;
        RECT 700.190 811.140 700.510 811.200 ;
        RECT 571.850 811.000 700.510 811.140 ;
        RECT 571.850 810.940 572.170 811.000 ;
        RECT 700.190 810.940 700.510 811.000 ;
      LAYER via ;
        RECT 700.220 3503.060 700.480 3503.320 ;
        RECT 770.600 3503.060 770.860 3503.320 ;
        RECT 571.880 810.940 572.140 811.200 ;
        RECT 700.220 810.940 700.480 811.200 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3503.350 770.800 3517.600 ;
        RECT 700.220 3503.030 700.480 3503.350 ;
        RECT 770.600 3503.030 770.860 3503.350 ;
        RECT 700.280 811.230 700.420 3503.030 ;
        RECT 571.880 810.910 572.140 811.230 ;
        RECT 700.220 810.910 700.480 811.230 ;
        RECT 570.290 799.410 570.570 800.000 ;
        RECT 571.940 799.410 572.080 810.910 ;
        RECT 570.290 799.270 572.080 799.410 ;
        RECT 570.290 796.000 570.570 799.270 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 441.670 832.560 441.990 832.620 ;
        RECT 575.530 832.560 575.850 832.620 ;
        RECT 441.670 832.420 575.850 832.560 ;
        RECT 441.670 832.360 441.990 832.420 ;
        RECT 575.530 832.360 575.850 832.420 ;
      LAYER via ;
        RECT 441.700 832.360 441.960 832.620 ;
        RECT 575.560 832.360 575.820 832.620 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3512.170 446.040 3517.600 ;
        RECT 441.760 3512.030 446.040 3512.170 ;
        RECT 441.760 832.650 441.900 3512.030 ;
        RECT 441.700 832.330 441.960 832.650 ;
        RECT 575.560 832.330 575.820 832.650 ;
        RECT 575.620 799.410 575.760 832.330 ;
        RECT 577.190 799.410 577.470 800.000 ;
        RECT 575.620 799.270 577.470 799.410 ;
        RECT 577.190 796.000 577.470 799.270 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 121.510 3502.240 121.830 3502.300 ;
        RECT 580.590 3502.240 580.910 3502.300 ;
        RECT 121.510 3502.100 580.910 3502.240 ;
        RECT 121.510 3502.040 121.830 3502.100 ;
        RECT 580.590 3502.040 580.910 3502.100 ;
      LAYER via ;
        RECT 121.540 3502.040 121.800 3502.300 ;
        RECT 580.620 3502.040 580.880 3502.300 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3502.330 121.740 3517.600 ;
        RECT 121.540 3502.010 121.800 3502.330 ;
        RECT 580.620 3502.010 580.880 3502.330 ;
        RECT 580.680 855.670 580.820 3502.010 ;
        RECT 580.680 855.530 582.660 855.670 ;
        RECT 582.520 799.410 582.660 855.530 ;
        RECT 584.090 799.410 584.370 800.000 ;
        RECT 582.520 799.270 584.370 799.410 ;
        RECT 584.090 796.000 584.370 799.270 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3354.000 17.410 3354.060 ;
        RECT 587.030 3354.000 587.350 3354.060 ;
        RECT 17.090 3353.860 587.350 3354.000 ;
        RECT 17.090 3353.800 17.410 3353.860 ;
        RECT 587.030 3353.800 587.350 3353.860 ;
        RECT 587.030 831.200 587.350 831.260 ;
        RECT 589.330 831.200 589.650 831.260 ;
        RECT 587.030 831.060 589.650 831.200 ;
        RECT 587.030 831.000 587.350 831.060 ;
        RECT 589.330 831.000 589.650 831.060 ;
      LAYER via ;
        RECT 17.120 3353.800 17.380 3354.060 ;
        RECT 587.060 3353.800 587.320 3354.060 ;
        RECT 587.060 831.000 587.320 831.260 ;
        RECT 589.360 831.000 589.620 831.260 ;
      LAYER met2 ;
        RECT 17.110 3355.955 17.390 3356.325 ;
        RECT 17.180 3354.090 17.320 3355.955 ;
        RECT 17.120 3353.770 17.380 3354.090 ;
        RECT 587.060 3353.770 587.320 3354.090 ;
        RECT 587.120 831.290 587.260 3353.770 ;
        RECT 587.060 830.970 587.320 831.290 ;
        RECT 589.360 830.970 589.620 831.290 ;
        RECT 589.420 799.410 589.560 830.970 ;
        RECT 590.990 799.410 591.270 800.000 ;
        RECT 589.420 799.270 591.270 799.410 ;
        RECT 590.990 796.000 591.270 799.270 ;
      LAYER via2 ;
        RECT 17.110 3356.000 17.390 3356.280 ;
      LAYER met3 ;
        RECT -4.800 3356.290 2.400 3356.740 ;
        RECT 17.085 3356.290 17.415 3356.305 ;
        RECT -4.800 3355.990 17.415 3356.290 ;
        RECT -4.800 3355.540 2.400 3355.990 ;
        RECT 17.085 3355.975 17.415 3355.990 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 3091.520 16.030 3091.580 ;
        RECT 589.790 3091.520 590.110 3091.580 ;
        RECT 15.710 3091.380 590.110 3091.520 ;
        RECT 15.710 3091.320 16.030 3091.380 ;
        RECT 589.790 3091.320 590.110 3091.380 ;
        RECT 589.790 821.000 590.110 821.060 ;
        RECT 596.230 821.000 596.550 821.060 ;
        RECT 589.790 820.860 596.550 821.000 ;
        RECT 589.790 820.800 590.110 820.860 ;
        RECT 596.230 820.800 596.550 820.860 ;
      LAYER via ;
        RECT 15.740 3091.320 16.000 3091.580 ;
        RECT 589.820 3091.320 590.080 3091.580 ;
        RECT 589.820 820.800 590.080 821.060 ;
        RECT 596.260 820.800 596.520 821.060 ;
      LAYER met2 ;
        RECT 15.730 3095.515 16.010 3095.885 ;
        RECT 15.800 3091.610 15.940 3095.515 ;
        RECT 15.740 3091.290 16.000 3091.610 ;
        RECT 589.820 3091.290 590.080 3091.610 ;
        RECT 589.880 821.090 590.020 3091.290 ;
        RECT 589.820 820.770 590.080 821.090 ;
        RECT 596.260 820.770 596.520 821.090 ;
        RECT 596.320 799.410 596.460 820.770 ;
        RECT 597.890 799.410 598.170 800.000 ;
        RECT 596.320 799.270 598.170 799.410 ;
        RECT 597.890 796.000 598.170 799.270 ;
      LAYER via2 ;
        RECT 15.730 3095.560 16.010 3095.840 ;
      LAYER met3 ;
        RECT -4.800 3095.850 2.400 3096.300 ;
        RECT 15.705 3095.850 16.035 3095.865 ;
        RECT -4.800 3095.550 16.035 3095.850 ;
        RECT -4.800 3095.100 2.400 3095.550 ;
        RECT 15.705 3095.535 16.035 3095.550 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2829.380 17.410 2829.440 ;
        RECT 600.830 2829.380 601.150 2829.440 ;
        RECT 17.090 2829.240 601.150 2829.380 ;
        RECT 17.090 2829.180 17.410 2829.240 ;
        RECT 600.830 2829.180 601.150 2829.240 ;
        RECT 600.830 815.900 601.150 815.960 ;
        RECT 603.130 815.900 603.450 815.960 ;
        RECT 600.830 815.760 603.450 815.900 ;
        RECT 600.830 815.700 601.150 815.760 ;
        RECT 603.130 815.700 603.450 815.760 ;
      LAYER via ;
        RECT 17.120 2829.180 17.380 2829.440 ;
        RECT 600.860 2829.180 601.120 2829.440 ;
        RECT 600.860 815.700 601.120 815.960 ;
        RECT 603.160 815.700 603.420 815.960 ;
      LAYER met2 ;
        RECT 17.110 2834.395 17.390 2834.765 ;
        RECT 17.180 2829.470 17.320 2834.395 ;
        RECT 17.120 2829.150 17.380 2829.470 ;
        RECT 600.860 2829.150 601.120 2829.470 ;
        RECT 600.920 815.990 601.060 2829.150 ;
        RECT 600.860 815.670 601.120 815.990 ;
        RECT 603.160 815.670 603.420 815.990 ;
        RECT 603.220 799.410 603.360 815.670 ;
        RECT 604.790 799.410 605.070 800.000 ;
        RECT 603.220 799.270 605.070 799.410 ;
        RECT 604.790 796.000 605.070 799.270 ;
      LAYER via2 ;
        RECT 17.110 2834.440 17.390 2834.720 ;
      LAYER met3 ;
        RECT -4.800 2834.730 2.400 2835.180 ;
        RECT 17.085 2834.730 17.415 2834.745 ;
        RECT -4.800 2834.430 17.415 2834.730 ;
        RECT -4.800 2833.980 2.400 2834.430 ;
        RECT 17.085 2834.415 17.415 2834.430 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2574.040 17.410 2574.100 ;
        RECT 607.730 2574.040 608.050 2574.100 ;
        RECT 17.090 2573.900 608.050 2574.040 ;
        RECT 17.090 2573.840 17.410 2573.900 ;
        RECT 607.730 2573.840 608.050 2573.900 ;
        RECT 607.730 815.900 608.050 815.960 ;
        RECT 610.030 815.900 610.350 815.960 ;
        RECT 607.730 815.760 610.350 815.900 ;
        RECT 607.730 815.700 608.050 815.760 ;
        RECT 610.030 815.700 610.350 815.760 ;
      LAYER via ;
        RECT 17.120 2573.840 17.380 2574.100 ;
        RECT 607.760 2573.840 608.020 2574.100 ;
        RECT 607.760 815.700 608.020 815.960 ;
        RECT 610.060 815.700 610.320 815.960 ;
      LAYER met2 ;
        RECT 17.110 2573.955 17.390 2574.325 ;
        RECT 17.120 2573.810 17.380 2573.955 ;
        RECT 607.760 2573.810 608.020 2574.130 ;
        RECT 607.820 815.990 607.960 2573.810 ;
        RECT 607.760 815.670 608.020 815.990 ;
        RECT 610.060 815.670 610.320 815.990 ;
        RECT 610.120 799.410 610.260 815.670 ;
        RECT 611.690 799.410 611.970 800.000 ;
        RECT 610.120 799.270 611.970 799.410 ;
        RECT 611.690 796.000 611.970 799.270 ;
      LAYER via2 ;
        RECT 17.110 2574.000 17.390 2574.280 ;
      LAYER met3 ;
        RECT -4.800 2574.290 2.400 2574.740 ;
        RECT 17.085 2574.290 17.415 2574.305 ;
        RECT -4.800 2573.990 17.415 2574.290 ;
        RECT -4.800 2573.540 2.400 2573.990 ;
        RECT 17.085 2573.975 17.415 2573.990 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 2311.900 16.490 2311.960 ;
        RECT 614.630 2311.900 614.950 2311.960 ;
        RECT 16.170 2311.760 614.950 2311.900 ;
        RECT 16.170 2311.700 16.490 2311.760 ;
        RECT 614.630 2311.700 614.950 2311.760 ;
        RECT 614.630 815.900 614.950 815.960 ;
        RECT 616.930 815.900 617.250 815.960 ;
        RECT 614.630 815.760 617.250 815.900 ;
        RECT 614.630 815.700 614.950 815.760 ;
        RECT 616.930 815.700 617.250 815.760 ;
      LAYER via ;
        RECT 16.200 2311.700 16.460 2311.960 ;
        RECT 614.660 2311.700 614.920 2311.960 ;
        RECT 614.660 815.700 614.920 815.960 ;
        RECT 616.960 815.700 617.220 815.960 ;
      LAYER met2 ;
        RECT 16.190 2312.835 16.470 2313.205 ;
        RECT 16.260 2311.990 16.400 2312.835 ;
        RECT 16.200 2311.670 16.460 2311.990 ;
        RECT 614.660 2311.670 614.920 2311.990 ;
        RECT 614.720 815.990 614.860 2311.670 ;
        RECT 614.660 815.670 614.920 815.990 ;
        RECT 616.960 815.670 617.220 815.990 ;
        RECT 617.020 799.410 617.160 815.670 ;
        RECT 618.590 799.410 618.870 800.000 ;
        RECT 617.020 799.270 618.870 799.410 ;
        RECT 618.590 796.000 618.870 799.270 ;
      LAYER via2 ;
        RECT 16.190 2312.880 16.470 2313.160 ;
      LAYER met3 ;
        RECT -4.800 2313.170 2.400 2313.620 ;
        RECT 16.165 2313.170 16.495 2313.185 ;
        RECT -4.800 2312.870 16.495 2313.170 ;
        RECT -4.800 2312.420 2.400 2312.870 ;
        RECT 16.165 2312.855 16.495 2312.870 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2049.420 16.030 2049.480 ;
        RECT 621.530 2049.420 621.850 2049.480 ;
        RECT 15.710 2049.280 621.850 2049.420 ;
        RECT 15.710 2049.220 16.030 2049.280 ;
        RECT 621.530 2049.220 621.850 2049.280 ;
        RECT 621.530 815.900 621.850 815.960 ;
        RECT 623.830 815.900 624.150 815.960 ;
        RECT 621.530 815.760 624.150 815.900 ;
        RECT 621.530 815.700 621.850 815.760 ;
        RECT 623.830 815.700 624.150 815.760 ;
      LAYER via ;
        RECT 15.740 2049.220 16.000 2049.480 ;
        RECT 621.560 2049.220 621.820 2049.480 ;
        RECT 621.560 815.700 621.820 815.960 ;
        RECT 623.860 815.700 624.120 815.960 ;
      LAYER met2 ;
        RECT 15.730 2052.395 16.010 2052.765 ;
        RECT 15.800 2049.510 15.940 2052.395 ;
        RECT 15.740 2049.190 16.000 2049.510 ;
        RECT 621.560 2049.190 621.820 2049.510 ;
        RECT 621.620 815.990 621.760 2049.190 ;
        RECT 621.560 815.670 621.820 815.990 ;
        RECT 623.860 815.670 624.120 815.990 ;
        RECT 623.920 799.410 624.060 815.670 ;
        RECT 625.490 799.410 625.770 800.000 ;
        RECT 623.920 799.270 625.770 799.410 ;
        RECT 625.490 796.000 625.770 799.270 ;
      LAYER via2 ;
        RECT 15.730 2052.440 16.010 2052.720 ;
      LAYER met3 ;
        RECT -4.800 2052.730 2.400 2053.180 ;
        RECT 15.705 2052.730 16.035 2052.745 ;
        RECT -4.800 2052.430 16.035 2052.730 ;
        RECT -4.800 2051.980 2.400 2052.430 ;
        RECT 15.705 2052.415 16.035 2052.430 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 439.830 796.660 440.150 796.920 ;
        RECT 439.920 794.140 440.060 796.660 ;
        RECT 686.850 794.140 687.170 794.200 ;
        RECT 439.920 794.000 687.170 794.140 ;
        RECT 686.850 793.940 687.170 794.000 ;
        RECT 686.850 503.440 687.170 503.500 ;
        RECT 2898.070 503.440 2898.390 503.500 ;
        RECT 686.850 503.300 2898.390 503.440 ;
        RECT 686.850 503.240 687.170 503.300 ;
        RECT 2898.070 503.240 2898.390 503.300 ;
      LAYER via ;
        RECT 439.860 796.660 440.120 796.920 ;
        RECT 686.880 793.940 687.140 794.200 ;
        RECT 686.880 503.240 687.140 503.500 ;
        RECT 2898.100 503.240 2898.360 503.500 ;
      LAYER met2 ;
        RECT 439.190 796.690 439.470 800.000 ;
        RECT 439.860 796.690 440.120 796.950 ;
        RECT 439.190 796.630 440.120 796.690 ;
        RECT 439.190 796.550 440.060 796.630 ;
        RECT 439.190 796.000 439.470 796.550 ;
        RECT 686.880 793.910 687.140 794.230 ;
        RECT 686.940 503.530 687.080 793.910 ;
        RECT 686.880 503.210 687.140 503.530 ;
        RECT 2898.100 503.210 2898.360 503.530 ;
        RECT 2898.160 497.605 2898.300 503.210 ;
        RECT 2898.090 497.235 2898.370 497.605 ;
      LAYER via2 ;
        RECT 2898.090 497.280 2898.370 497.560 ;
      LAYER met3 ;
        RECT 2898.065 497.570 2898.395 497.585 ;
        RECT 2917.600 497.570 2924.800 498.020 ;
        RECT 2898.065 497.270 2924.800 497.570 ;
        RECT 2898.065 497.255 2898.395 497.270 ;
        RECT 2917.600 496.820 2924.800 497.270 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 1787.280 16.030 1787.340 ;
        RECT 628.430 1787.280 628.750 1787.340 ;
        RECT 15.710 1787.140 628.750 1787.280 ;
        RECT 15.710 1787.080 16.030 1787.140 ;
        RECT 628.430 1787.080 628.750 1787.140 ;
        RECT 628.430 815.900 628.750 815.960 ;
        RECT 630.730 815.900 631.050 815.960 ;
        RECT 628.430 815.760 631.050 815.900 ;
        RECT 628.430 815.700 628.750 815.760 ;
        RECT 630.730 815.700 631.050 815.760 ;
      LAYER via ;
        RECT 15.740 1787.080 16.000 1787.340 ;
        RECT 628.460 1787.080 628.720 1787.340 ;
        RECT 628.460 815.700 628.720 815.960 ;
        RECT 630.760 815.700 631.020 815.960 ;
      LAYER met2 ;
        RECT 15.730 1791.955 16.010 1792.325 ;
        RECT 15.800 1787.370 15.940 1791.955 ;
        RECT 15.740 1787.050 16.000 1787.370 ;
        RECT 628.460 1787.050 628.720 1787.370 ;
        RECT 628.520 815.990 628.660 1787.050 ;
        RECT 628.460 815.670 628.720 815.990 ;
        RECT 630.760 815.670 631.020 815.990 ;
        RECT 630.820 799.410 630.960 815.670 ;
        RECT 632.390 799.410 632.670 800.000 ;
        RECT 630.820 799.270 632.670 799.410 ;
        RECT 632.390 796.000 632.670 799.270 ;
      LAYER via2 ;
        RECT 15.730 1792.000 16.010 1792.280 ;
      LAYER met3 ;
        RECT -4.800 1792.290 2.400 1792.740 ;
        RECT 15.705 1792.290 16.035 1792.305 ;
        RECT -4.800 1791.990 16.035 1792.290 ;
        RECT -4.800 1791.540 2.400 1791.990 ;
        RECT 15.705 1791.975 16.035 1791.990 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 1525.140 16.490 1525.200 ;
        RECT 635.330 1525.140 635.650 1525.200 ;
        RECT 16.170 1525.000 635.650 1525.140 ;
        RECT 16.170 1524.940 16.490 1525.000 ;
        RECT 635.330 1524.940 635.650 1525.000 ;
        RECT 635.330 815.900 635.650 815.960 ;
        RECT 637.630 815.900 637.950 815.960 ;
        RECT 635.330 815.760 637.950 815.900 ;
        RECT 635.330 815.700 635.650 815.760 ;
        RECT 637.630 815.700 637.950 815.760 ;
      LAYER via ;
        RECT 16.200 1524.940 16.460 1525.200 ;
        RECT 635.360 1524.940 635.620 1525.200 ;
        RECT 635.360 815.700 635.620 815.960 ;
        RECT 637.660 815.700 637.920 815.960 ;
      LAYER met2 ;
        RECT 16.190 1530.835 16.470 1531.205 ;
        RECT 16.260 1525.230 16.400 1530.835 ;
        RECT 16.200 1524.910 16.460 1525.230 ;
        RECT 635.360 1524.910 635.620 1525.230 ;
        RECT 635.420 815.990 635.560 1524.910 ;
        RECT 635.360 815.670 635.620 815.990 ;
        RECT 637.660 815.670 637.920 815.990 ;
        RECT 637.720 799.410 637.860 815.670 ;
        RECT 639.290 799.410 639.570 800.000 ;
        RECT 637.720 799.270 639.570 799.410 ;
        RECT 639.290 796.000 639.570 799.270 ;
      LAYER via2 ;
        RECT 16.190 1530.880 16.470 1531.160 ;
      LAYER met3 ;
        RECT -4.800 1531.170 2.400 1531.620 ;
        RECT 16.165 1531.170 16.495 1531.185 ;
        RECT -4.800 1530.870 16.495 1531.170 ;
        RECT -4.800 1530.420 2.400 1530.870 ;
        RECT 16.165 1530.855 16.495 1530.870 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 1269.800 17.410 1269.860 ;
        RECT 642.230 1269.800 642.550 1269.860 ;
        RECT 17.090 1269.660 642.550 1269.800 ;
        RECT 17.090 1269.600 17.410 1269.660 ;
        RECT 642.230 1269.600 642.550 1269.660 ;
        RECT 642.230 831.200 642.550 831.260 ;
        RECT 644.530 831.200 644.850 831.260 ;
        RECT 642.230 831.060 644.850 831.200 ;
        RECT 642.230 831.000 642.550 831.060 ;
        RECT 644.530 831.000 644.850 831.060 ;
      LAYER via ;
        RECT 17.120 1269.600 17.380 1269.860 ;
        RECT 642.260 1269.600 642.520 1269.860 ;
        RECT 642.260 831.000 642.520 831.260 ;
        RECT 644.560 831.000 644.820 831.260 ;
      LAYER met2 ;
        RECT 17.110 1270.395 17.390 1270.765 ;
        RECT 17.180 1269.890 17.320 1270.395 ;
        RECT 17.120 1269.570 17.380 1269.890 ;
        RECT 642.260 1269.570 642.520 1269.890 ;
        RECT 642.320 831.290 642.460 1269.570 ;
        RECT 642.260 830.970 642.520 831.290 ;
        RECT 644.560 830.970 644.820 831.290 ;
        RECT 644.620 799.410 644.760 830.970 ;
        RECT 646.190 799.410 646.470 800.000 ;
        RECT 644.620 799.270 646.470 799.410 ;
        RECT 646.190 796.000 646.470 799.270 ;
      LAYER via2 ;
        RECT 17.110 1270.440 17.390 1270.720 ;
      LAYER met3 ;
        RECT -4.800 1270.730 2.400 1271.180 ;
        RECT 17.085 1270.730 17.415 1270.745 ;
        RECT -4.800 1270.430 17.415 1270.730 ;
        RECT -4.800 1269.980 2.400 1270.430 ;
        RECT 17.085 1270.415 17.415 1270.430 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 1007.660 17.410 1007.720 ;
        RECT 649.130 1007.660 649.450 1007.720 ;
        RECT 17.090 1007.520 649.450 1007.660 ;
        RECT 17.090 1007.460 17.410 1007.520 ;
        RECT 649.130 1007.460 649.450 1007.520 ;
        RECT 649.130 831.200 649.450 831.260 ;
        RECT 651.430 831.200 651.750 831.260 ;
        RECT 649.130 831.060 651.750 831.200 ;
        RECT 649.130 831.000 649.450 831.060 ;
        RECT 651.430 831.000 651.750 831.060 ;
      LAYER via ;
        RECT 17.120 1007.460 17.380 1007.720 ;
        RECT 649.160 1007.460 649.420 1007.720 ;
        RECT 649.160 831.000 649.420 831.260 ;
        RECT 651.460 831.000 651.720 831.260 ;
      LAYER met2 ;
        RECT 17.110 1009.275 17.390 1009.645 ;
        RECT 17.180 1007.750 17.320 1009.275 ;
        RECT 17.120 1007.430 17.380 1007.750 ;
        RECT 649.160 1007.430 649.420 1007.750 ;
        RECT 649.220 831.290 649.360 1007.430 ;
        RECT 649.160 830.970 649.420 831.290 ;
        RECT 651.460 830.970 651.720 831.290 ;
        RECT 651.520 799.410 651.660 830.970 ;
        RECT 653.090 799.410 653.370 800.000 ;
        RECT 651.520 799.270 653.370 799.410 ;
        RECT 653.090 796.000 653.370 799.270 ;
      LAYER via2 ;
        RECT 17.110 1009.320 17.390 1009.600 ;
      LAYER met3 ;
        RECT -4.800 1009.610 2.400 1010.060 ;
        RECT 17.085 1009.610 17.415 1009.625 ;
        RECT -4.800 1009.310 17.415 1009.610 ;
        RECT -4.800 1008.860 2.400 1009.310 ;
        RECT 17.085 1009.295 17.415 1009.310 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 44.690 808.760 45.010 808.820 ;
        RECT 658.330 808.760 658.650 808.820 ;
        RECT 44.690 808.620 658.650 808.760 ;
        RECT 44.690 808.560 45.010 808.620 ;
        RECT 658.330 808.560 658.650 808.620 ;
        RECT 16.630 751.980 16.950 752.040 ;
        RECT 44.690 751.980 45.010 752.040 ;
        RECT 16.630 751.840 45.010 751.980 ;
        RECT 16.630 751.780 16.950 751.840 ;
        RECT 44.690 751.780 45.010 751.840 ;
      LAYER via ;
        RECT 44.720 808.560 44.980 808.820 ;
        RECT 658.360 808.560 658.620 808.820 ;
        RECT 16.660 751.780 16.920 752.040 ;
        RECT 44.720 751.780 44.980 752.040 ;
      LAYER met2 ;
        RECT 44.720 808.530 44.980 808.850 ;
        RECT 658.360 808.530 658.620 808.850 ;
        RECT 44.780 752.070 44.920 808.530 ;
        RECT 658.420 799.410 658.560 808.530 ;
        RECT 659.990 799.410 660.270 800.000 ;
        RECT 658.420 799.270 660.270 799.410 ;
        RECT 659.990 796.000 660.270 799.270 ;
        RECT 16.660 751.750 16.920 752.070 ;
        RECT 44.720 751.750 44.980 752.070 ;
        RECT 16.720 749.205 16.860 751.750 ;
        RECT 16.650 748.835 16.930 749.205 ;
      LAYER via2 ;
        RECT 16.650 748.880 16.930 749.160 ;
      LAYER met3 ;
        RECT -4.800 749.170 2.400 749.620 ;
        RECT 16.625 749.170 16.955 749.185 ;
        RECT -4.800 748.870 16.955 749.170 ;
        RECT -4.800 748.420 2.400 748.870 ;
        RECT 16.625 748.855 16.955 748.870 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 603.590 809.780 603.910 809.840 ;
        RECT 665.230 809.780 665.550 809.840 ;
        RECT 603.590 809.640 665.550 809.780 ;
        RECT 603.590 809.580 603.910 809.640 ;
        RECT 665.230 809.580 665.550 809.640 ;
        RECT 51.590 809.100 51.910 809.160 ;
        RECT 603.590 809.100 603.910 809.160 ;
        RECT 51.590 808.960 603.910 809.100 ;
        RECT 51.590 808.900 51.910 808.960 ;
        RECT 603.590 808.900 603.910 808.960 ;
        RECT 16.630 489.840 16.950 489.900 ;
        RECT 51.590 489.840 51.910 489.900 ;
        RECT 16.630 489.700 51.910 489.840 ;
        RECT 16.630 489.640 16.950 489.700 ;
        RECT 51.590 489.640 51.910 489.700 ;
      LAYER via ;
        RECT 603.620 809.580 603.880 809.840 ;
        RECT 665.260 809.580 665.520 809.840 ;
        RECT 51.620 808.900 51.880 809.160 ;
        RECT 603.620 808.900 603.880 809.160 ;
        RECT 16.660 489.640 16.920 489.900 ;
        RECT 51.620 489.640 51.880 489.900 ;
      LAYER met2 ;
        RECT 603.620 809.550 603.880 809.870 ;
        RECT 665.260 809.550 665.520 809.870 ;
        RECT 603.680 809.190 603.820 809.550 ;
        RECT 51.620 808.870 51.880 809.190 ;
        RECT 603.620 808.870 603.880 809.190 ;
        RECT 51.680 489.930 51.820 808.870 ;
        RECT 665.320 799.410 665.460 809.550 ;
        RECT 666.890 799.410 667.170 800.000 ;
        RECT 665.320 799.270 667.170 799.410 ;
        RECT 666.890 796.000 667.170 799.270 ;
        RECT 16.660 489.610 16.920 489.930 ;
        RECT 51.620 489.610 51.880 489.930 ;
        RECT 16.720 488.085 16.860 489.610 ;
        RECT 16.650 487.715 16.930 488.085 ;
      LAYER via2 ;
        RECT 16.650 487.760 16.930 488.040 ;
      LAYER met3 ;
        RECT -4.800 488.050 2.400 488.500 ;
        RECT 16.625 488.050 16.955 488.065 ;
        RECT -4.800 487.750 16.955 488.050 ;
        RECT -4.800 487.300 2.400 487.750 ;
        RECT 16.625 487.735 16.955 487.750 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 808.080 18.330 808.140 ;
        RECT 672.130 808.080 672.450 808.140 ;
        RECT 18.010 807.940 672.450 808.080 ;
        RECT 18.010 807.880 18.330 807.940 ;
        RECT 672.130 807.880 672.450 807.940 ;
      LAYER via ;
        RECT 18.040 807.880 18.300 808.140 ;
        RECT 672.160 807.880 672.420 808.140 ;
      LAYER met2 ;
        RECT 18.040 807.850 18.300 808.170 ;
        RECT 672.160 807.850 672.420 808.170 ;
        RECT 18.100 292.925 18.240 807.850 ;
        RECT 672.220 799.410 672.360 807.850 ;
        RECT 673.790 799.410 674.070 800.000 ;
        RECT 672.220 799.270 674.070 799.410 ;
        RECT 673.790 796.000 674.070 799.270 ;
        RECT 18.030 292.555 18.310 292.925 ;
      LAYER via2 ;
        RECT 18.030 292.600 18.310 292.880 ;
      LAYER met3 ;
        RECT -4.800 292.890 2.400 293.340 ;
        RECT 18.005 292.890 18.335 292.905 ;
        RECT -4.800 292.590 18.335 292.890 ;
        RECT -4.800 292.140 2.400 292.590 ;
        RECT 18.005 292.575 18.335 292.590 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 103.260 17.410 103.320 ;
        RECT 681.790 103.260 682.110 103.320 ;
        RECT 17.090 103.120 682.110 103.260 ;
        RECT 17.090 103.060 17.410 103.120 ;
        RECT 681.790 103.060 682.110 103.120 ;
      LAYER via ;
        RECT 17.120 103.060 17.380 103.320 ;
        RECT 681.820 103.060 682.080 103.320 ;
      LAYER met2 ;
        RECT 680.690 796.690 680.970 800.000 ;
        RECT 680.690 796.550 682.020 796.690 ;
        RECT 680.690 796.000 680.970 796.550 ;
        RECT 681.880 103.350 682.020 796.550 ;
        RECT 17.120 103.030 17.380 103.350 ;
        RECT 681.820 103.030 682.080 103.350 ;
        RECT 17.180 97.085 17.320 103.030 ;
        RECT 17.110 96.715 17.390 97.085 ;
      LAYER via2 ;
        RECT 17.110 96.760 17.390 97.040 ;
      LAYER met3 ;
        RECT -4.800 97.050 2.400 97.500 ;
        RECT 17.085 97.050 17.415 97.065 ;
        RECT -4.800 96.750 17.415 97.050 ;
        RECT -4.800 96.300 2.400 96.750 ;
        RECT 17.085 96.735 17.415 96.750 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 447.190 809.440 447.510 809.500 ;
        RECT 693.750 809.440 694.070 809.500 ;
        RECT 447.190 809.300 604.280 809.440 ;
        RECT 447.190 809.240 447.510 809.300 ;
        RECT 604.140 809.100 604.280 809.300 ;
        RECT 627.830 809.300 694.070 809.440 ;
        RECT 627.830 809.100 627.970 809.300 ;
        RECT 693.750 809.240 694.070 809.300 ;
        RECT 604.140 808.960 627.970 809.100 ;
        RECT 695.130 696.900 695.450 696.960 ;
        RECT 2900.830 696.900 2901.150 696.960 ;
        RECT 695.130 696.760 2901.150 696.900 ;
        RECT 695.130 696.700 695.450 696.760 ;
        RECT 2900.830 696.700 2901.150 696.760 ;
      LAYER via ;
        RECT 447.220 809.240 447.480 809.500 ;
        RECT 693.780 809.240 694.040 809.500 ;
        RECT 695.160 696.700 695.420 696.960 ;
        RECT 2900.860 696.700 2901.120 696.960 ;
      LAYER met2 ;
        RECT 447.220 809.210 447.480 809.530 ;
        RECT 693.780 809.210 694.040 809.530 ;
        RECT 446.090 799.410 446.370 800.000 ;
        RECT 447.280 799.410 447.420 809.210 ;
        RECT 446.090 799.270 447.420 799.410 ;
        RECT 446.090 796.000 446.370 799.270 ;
        RECT 693.840 759.070 693.980 809.210 ;
        RECT 693.840 758.930 695.360 759.070 ;
        RECT 695.220 696.990 695.360 758.930 ;
        RECT 695.160 696.670 695.420 696.990 ;
        RECT 2900.860 696.845 2901.120 696.990 ;
        RECT 2900.850 696.475 2901.130 696.845 ;
      LAYER via2 ;
        RECT 2900.850 696.520 2901.130 696.800 ;
      LAYER met3 ;
        RECT 2900.825 696.810 2901.155 696.825 ;
        RECT 2917.600 696.810 2924.800 697.260 ;
        RECT 2900.825 696.510 2924.800 696.810 ;
        RECT 2900.825 696.495 2901.155 696.510 ;
        RECT 2917.600 696.060 2924.800 696.510 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 449.490 890.360 449.810 890.420 ;
        RECT 2900.830 890.360 2901.150 890.420 ;
        RECT 449.490 890.220 2901.150 890.360 ;
        RECT 449.490 890.160 449.810 890.220 ;
        RECT 2900.830 890.160 2901.150 890.220 ;
      LAYER via ;
        RECT 449.520 890.160 449.780 890.420 ;
        RECT 2900.860 890.160 2901.120 890.420 ;
      LAYER met2 ;
        RECT 2900.850 895.715 2901.130 896.085 ;
        RECT 2900.920 890.450 2901.060 895.715 ;
        RECT 449.520 890.130 449.780 890.450 ;
        RECT 2900.860 890.130 2901.120 890.450 ;
        RECT 449.580 855.670 449.720 890.130 ;
        RECT 449.580 855.530 451.560 855.670 ;
        RECT 451.420 799.410 451.560 855.530 ;
        RECT 452.990 799.410 453.270 800.000 ;
        RECT 451.420 799.270 453.270 799.410 ;
        RECT 452.990 796.000 453.270 799.270 ;
      LAYER via2 ;
        RECT 2900.850 895.760 2901.130 896.040 ;
      LAYER met3 ;
        RECT 2900.825 896.050 2901.155 896.065 ;
        RECT 2917.600 896.050 2924.800 896.500 ;
        RECT 2900.825 895.750 2924.800 896.050 ;
        RECT 2900.825 895.735 2901.155 895.750 ;
        RECT 2917.600 895.300 2924.800 895.750 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.390 1090.280 456.710 1090.340 ;
        RECT 2900.830 1090.280 2901.150 1090.340 ;
        RECT 456.390 1090.140 2901.150 1090.280 ;
        RECT 456.390 1090.080 456.710 1090.140 ;
        RECT 2900.830 1090.080 2901.150 1090.140 ;
      LAYER via ;
        RECT 456.420 1090.080 456.680 1090.340 ;
        RECT 2900.860 1090.080 2901.120 1090.340 ;
      LAYER met2 ;
        RECT 2900.850 1094.955 2901.130 1095.325 ;
        RECT 2900.920 1090.370 2901.060 1094.955 ;
        RECT 456.420 1090.050 456.680 1090.370 ;
        RECT 2900.860 1090.050 2901.120 1090.370 ;
        RECT 456.480 855.670 456.620 1090.050 ;
        RECT 456.480 855.530 458.460 855.670 ;
        RECT 458.320 799.410 458.460 855.530 ;
        RECT 459.890 799.410 460.170 800.000 ;
        RECT 458.320 799.270 460.170 799.410 ;
        RECT 459.890 796.000 460.170 799.270 ;
      LAYER via2 ;
        RECT 2900.850 1095.000 2901.130 1095.280 ;
      LAYER met3 ;
        RECT 2900.825 1095.290 2901.155 1095.305 ;
        RECT 2917.600 1095.290 2924.800 1095.740 ;
        RECT 2900.825 1094.990 2924.800 1095.290 ;
        RECT 2900.825 1094.975 2901.155 1094.990 ;
        RECT 2917.600 1094.540 2924.800 1094.990 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 463.290 1290.540 463.610 1290.600 ;
        RECT 2900.830 1290.540 2901.150 1290.600 ;
        RECT 463.290 1290.400 2901.150 1290.540 ;
        RECT 463.290 1290.340 463.610 1290.400 ;
        RECT 2900.830 1290.340 2901.150 1290.400 ;
      LAYER via ;
        RECT 463.320 1290.340 463.580 1290.600 ;
        RECT 2900.860 1290.340 2901.120 1290.600 ;
      LAYER met2 ;
        RECT 2900.850 1294.195 2901.130 1294.565 ;
        RECT 2900.920 1290.630 2901.060 1294.195 ;
        RECT 463.320 1290.310 463.580 1290.630 ;
        RECT 2900.860 1290.310 2901.120 1290.630 ;
        RECT 463.380 855.670 463.520 1290.310 ;
        RECT 463.380 855.530 465.360 855.670 ;
        RECT 465.220 799.410 465.360 855.530 ;
        RECT 466.790 799.410 467.070 800.000 ;
        RECT 465.220 799.270 467.070 799.410 ;
        RECT 466.790 796.000 467.070 799.270 ;
      LAYER via2 ;
        RECT 2900.850 1294.240 2901.130 1294.520 ;
      LAYER met3 ;
        RECT 2900.825 1294.530 2901.155 1294.545 ;
        RECT 2917.600 1294.530 2924.800 1294.980 ;
        RECT 2900.825 1294.230 2924.800 1294.530 ;
        RECT 2900.825 1294.215 2901.155 1294.230 ;
        RECT 2917.600 1293.780 2924.800 1294.230 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 470.190 1559.480 470.510 1559.540 ;
        RECT 2900.830 1559.480 2901.150 1559.540 ;
        RECT 470.190 1559.340 2901.150 1559.480 ;
        RECT 470.190 1559.280 470.510 1559.340 ;
        RECT 2900.830 1559.280 2901.150 1559.340 ;
      LAYER via ;
        RECT 470.220 1559.280 470.480 1559.540 ;
        RECT 2900.860 1559.280 2901.120 1559.540 ;
      LAYER met2 ;
        RECT 2900.850 1560.075 2901.130 1560.445 ;
        RECT 2900.920 1559.570 2901.060 1560.075 ;
        RECT 470.220 1559.250 470.480 1559.570 ;
        RECT 2900.860 1559.250 2901.120 1559.570 ;
        RECT 470.280 855.670 470.420 1559.250 ;
        RECT 470.280 855.530 472.260 855.670 ;
        RECT 472.120 799.410 472.260 855.530 ;
        RECT 473.690 799.410 473.970 800.000 ;
        RECT 472.120 799.270 473.970 799.410 ;
        RECT 473.690 796.000 473.970 799.270 ;
      LAYER via2 ;
        RECT 2900.850 1560.120 2901.130 1560.400 ;
      LAYER met3 ;
        RECT 2900.825 1560.410 2901.155 1560.425 ;
        RECT 2917.600 1560.410 2924.800 1560.860 ;
        RECT 2900.825 1560.110 2924.800 1560.410 ;
        RECT 2900.825 1560.095 2901.155 1560.110 ;
        RECT 2917.600 1559.660 2924.800 1560.110 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 477.090 1821.960 477.410 1822.020 ;
        RECT 2900.830 1821.960 2901.150 1822.020 ;
        RECT 477.090 1821.820 2901.150 1821.960 ;
        RECT 477.090 1821.760 477.410 1821.820 ;
        RECT 2900.830 1821.760 2901.150 1821.820 ;
      LAYER via ;
        RECT 477.120 1821.760 477.380 1822.020 ;
        RECT 2900.860 1821.760 2901.120 1822.020 ;
      LAYER met2 ;
        RECT 2900.850 1825.275 2901.130 1825.645 ;
        RECT 2900.920 1822.050 2901.060 1825.275 ;
        RECT 477.120 1821.730 477.380 1822.050 ;
        RECT 2900.860 1821.730 2901.120 1822.050 ;
        RECT 477.180 855.670 477.320 1821.730 ;
        RECT 477.180 855.530 479.160 855.670 ;
        RECT 479.020 799.410 479.160 855.530 ;
        RECT 480.590 799.410 480.870 800.000 ;
        RECT 479.020 799.270 480.870 799.410 ;
        RECT 480.590 796.000 480.870 799.270 ;
      LAYER via2 ;
        RECT 2900.850 1825.320 2901.130 1825.600 ;
      LAYER met3 ;
        RECT 2900.825 1825.610 2901.155 1825.625 ;
        RECT 2917.600 1825.610 2924.800 1826.060 ;
        RECT 2900.825 1825.310 2924.800 1825.610 ;
        RECT 2900.825 1825.295 2901.155 1825.310 ;
        RECT 2917.600 1824.860 2924.800 1825.310 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.990 2090.900 484.310 2090.960 ;
        RECT 2900.830 2090.900 2901.150 2090.960 ;
        RECT 483.990 2090.760 2901.150 2090.900 ;
        RECT 483.990 2090.700 484.310 2090.760 ;
        RECT 2900.830 2090.700 2901.150 2090.760 ;
      LAYER via ;
        RECT 484.020 2090.700 484.280 2090.960 ;
        RECT 2900.860 2090.700 2901.120 2090.960 ;
      LAYER met2 ;
        RECT 2900.850 2091.155 2901.130 2091.525 ;
        RECT 2900.920 2090.990 2901.060 2091.155 ;
        RECT 484.020 2090.670 484.280 2090.990 ;
        RECT 2900.860 2090.670 2901.120 2090.990 ;
        RECT 484.080 855.670 484.220 2090.670 ;
        RECT 484.080 855.530 486.060 855.670 ;
        RECT 485.920 799.410 486.060 855.530 ;
        RECT 487.490 799.410 487.770 800.000 ;
        RECT 485.920 799.270 487.770 799.410 ;
        RECT 487.490 796.000 487.770 799.270 ;
      LAYER via2 ;
        RECT 2900.850 2091.200 2901.130 2091.480 ;
      LAYER met3 ;
        RECT 2900.825 2091.490 2901.155 2091.505 ;
        RECT 2917.600 2091.490 2924.800 2091.940 ;
        RECT 2900.825 2091.190 2924.800 2091.490 ;
        RECT 2900.825 2091.175 2901.155 2091.190 ;
        RECT 2917.600 2090.740 2924.800 2091.190 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 485.140 499.500 485.460 499.760 ;
        RECT 485.230 498.680 485.370 499.500 ;
        RECT 485.230 498.540 486.520 498.680 ;
        RECT 483.990 497.320 484.310 497.380 ;
        RECT 486.380 497.320 486.520 498.540 ;
        RECT 483.990 497.180 486.520 497.320 ;
        RECT 483.990 497.120 484.310 497.180 ;
        RECT 629.350 19.960 629.670 20.020 ;
        RECT 524.560 19.820 629.670 19.960 ;
        RECT 483.990 19.620 484.310 19.680 ;
        RECT 524.560 19.620 524.700 19.820 ;
        RECT 629.350 19.760 629.670 19.820 ;
        RECT 483.990 19.480 524.700 19.620 ;
        RECT 483.990 19.420 484.310 19.480 ;
      LAYER via ;
        RECT 485.170 499.500 485.430 499.760 ;
        RECT 484.020 497.120 484.280 497.380 ;
        RECT 484.020 19.420 484.280 19.680 ;
        RECT 629.380 19.760 629.640 20.020 ;
      LAYER met2 ;
        RECT 485.190 500.000 485.470 504.000 ;
        RECT 485.230 499.790 485.370 500.000 ;
        RECT 485.170 499.470 485.430 499.790 ;
        RECT 484.020 497.090 484.280 497.410 ;
        RECT 484.080 19.710 484.220 497.090 ;
        RECT 629.380 19.730 629.640 20.050 ;
        RECT 484.020 19.390 484.280 19.710 ;
        RECT 629.440 2.400 629.580 19.730 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.190 500.000 623.470 504.000 ;
        RECT 623.230 499.645 623.370 500.000 ;
        RECT 623.160 499.275 623.440 499.645 ;
        RECT 2401.290 486.355 2401.570 486.725 ;
        RECT 2401.360 82.870 2401.500 486.355 ;
        RECT 2401.360 82.730 2402.880 82.870 ;
        RECT 2402.740 2.400 2402.880 82.730 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
      LAYER via2 ;
        RECT 623.160 499.320 623.440 499.600 ;
        RECT 2401.290 486.400 2401.570 486.680 ;
      LAYER met3 ;
        RECT 623.135 499.620 623.465 499.625 ;
        RECT 623.110 499.610 623.490 499.620 ;
        RECT 623.110 499.310 623.920 499.610 ;
        RECT 623.110 499.300 623.490 499.310 ;
        RECT 623.135 499.295 623.465 499.300 ;
        RECT 623.110 486.690 623.490 486.700 ;
        RECT 2401.265 486.690 2401.595 486.705 ;
        RECT 623.110 486.390 2401.595 486.690 ;
        RECT 623.110 486.380 623.490 486.390 ;
        RECT 2401.265 486.375 2401.595 486.390 ;
      LAYER via3 ;
        RECT 623.140 499.300 623.460 499.620 ;
        RECT 623.140 486.380 623.460 486.700 ;
      LAYER met4 ;
        RECT 623.135 499.295 623.465 499.625 ;
        RECT 623.150 486.705 623.450 499.295 ;
        RECT 623.135 486.375 623.465 486.705 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.070 472.840 621.390 472.900 ;
        RECT 623.370 472.840 623.690 472.900 ;
        RECT 621.070 472.700 623.690 472.840 ;
        RECT 621.070 472.640 621.390 472.700 ;
        RECT 623.370 472.640 623.690 472.700 ;
        RECT 621.070 17.920 621.390 17.980 ;
        RECT 2420.130 17.920 2420.450 17.980 ;
        RECT 621.070 17.780 2420.450 17.920 ;
        RECT 621.070 17.720 621.390 17.780 ;
        RECT 2420.130 17.720 2420.450 17.780 ;
      LAYER via ;
        RECT 621.100 472.640 621.360 472.900 ;
        RECT 623.400 472.640 623.660 472.900 ;
        RECT 621.100 17.720 621.360 17.980 ;
        RECT 2420.160 17.720 2420.420 17.980 ;
      LAYER met2 ;
        RECT 624.570 500.000 624.850 504.000 ;
        RECT 624.610 498.680 624.750 500.000 ;
        RECT 623.460 498.540 624.750 498.680 ;
        RECT 623.460 472.930 623.600 498.540 ;
        RECT 621.100 472.610 621.360 472.930 ;
        RECT 623.400 472.610 623.660 472.930 ;
        RECT 621.160 18.010 621.300 472.610 ;
        RECT 621.100 17.690 621.360 18.010 ;
        RECT 2420.160 17.690 2420.420 18.010 ;
        RECT 2420.220 2.400 2420.360 17.690 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.950 500.000 626.230 504.000 ;
        RECT 625.990 499.645 626.130 500.000 ;
        RECT 625.920 499.275 626.200 499.645 ;
        RECT 2438.090 17.835 2438.370 18.205 ;
        RECT 2438.160 2.400 2438.300 17.835 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
      LAYER via2 ;
        RECT 625.920 499.320 626.200 499.600 ;
        RECT 2438.090 17.880 2438.370 18.160 ;
      LAYER met3 ;
        RECT 625.895 499.620 626.225 499.625 ;
        RECT 625.870 499.610 626.250 499.620 ;
        RECT 625.440 499.310 626.250 499.610 ;
        RECT 625.870 499.300 626.250 499.310 ;
        RECT 625.895 499.295 626.225 499.300 ;
        RECT 625.870 18.170 626.250 18.180 ;
        RECT 2438.065 18.170 2438.395 18.185 ;
        RECT 625.870 17.870 2438.395 18.170 ;
        RECT 625.870 17.860 626.250 17.870 ;
        RECT 2438.065 17.855 2438.395 17.870 ;
      LAYER via3 ;
        RECT 625.900 499.300 626.220 499.620 ;
        RECT 625.900 17.860 626.220 18.180 ;
      LAYER met4 ;
        RECT 625.895 499.295 626.225 499.625 ;
        RECT 625.910 18.185 626.210 499.295 ;
        RECT 625.895 17.855 626.225 18.185 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.330 500.000 627.610 504.000 ;
        RECT 627.370 498.680 627.510 500.000 ;
        RECT 627.140 498.540 627.510 498.680 ;
        RECT 627.140 483.325 627.280 498.540 ;
        RECT 627.070 482.955 627.350 483.325 ;
        RECT 2455.570 17.155 2455.850 17.525 ;
        RECT 2455.640 2.400 2455.780 17.155 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
      LAYER via2 ;
        RECT 627.070 483.000 627.350 483.280 ;
        RECT 2455.570 17.200 2455.850 17.480 ;
      LAYER met3 ;
        RECT 627.045 483.300 627.375 483.305 ;
        RECT 626.790 483.290 627.375 483.300 ;
        RECT 626.590 482.990 627.375 483.290 ;
        RECT 626.790 482.980 627.375 482.990 ;
        RECT 627.045 482.975 627.375 482.980 ;
        RECT 626.790 17.490 627.170 17.500 ;
        RECT 2455.545 17.490 2455.875 17.505 ;
        RECT 626.790 17.190 2455.875 17.490 ;
        RECT 626.790 17.180 627.170 17.190 ;
        RECT 2455.545 17.175 2455.875 17.190 ;
      LAYER via3 ;
        RECT 626.820 482.980 627.140 483.300 ;
        RECT 626.820 17.180 627.140 17.500 ;
      LAYER met4 ;
        RECT 626.815 482.975 627.145 483.305 ;
        RECT 626.830 17.505 627.130 482.975 ;
        RECT 626.815 17.175 627.145 17.505 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 627.510 487.800 627.830 487.860 ;
        RECT 627.510 487.660 665.920 487.800 ;
        RECT 627.510 487.600 627.830 487.660 ;
        RECT 665.780 487.120 665.920 487.660 ;
        RECT 2470.270 487.120 2470.590 487.180 ;
        RECT 665.780 486.980 2470.590 487.120 ;
        RECT 2470.270 486.920 2470.590 486.980 ;
      LAYER via ;
        RECT 627.540 487.600 627.800 487.860 ;
        RECT 2470.300 486.920 2470.560 487.180 ;
      LAYER met2 ;
        RECT 628.710 500.000 628.990 504.000 ;
        RECT 628.750 498.850 628.890 500.000 ;
        RECT 628.520 498.710 628.890 498.850 ;
        RECT 628.520 498.000 628.660 498.710 ;
        RECT 627.830 497.860 628.660 498.000 ;
        RECT 627.830 497.490 627.970 497.860 ;
        RECT 627.600 497.350 627.970 497.490 ;
        RECT 627.600 487.890 627.740 497.350 ;
        RECT 627.540 487.570 627.800 487.890 ;
        RECT 2470.300 486.890 2470.560 487.210 ;
        RECT 2470.360 82.870 2470.500 486.890 ;
        RECT 2470.360 82.730 2473.720 82.870 ;
        RECT 2473.580 2.400 2473.720 82.730 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 630.040 499.700 630.360 499.760 ;
        RECT 629.210 499.560 630.360 499.700 ;
        RECT 629.210 498.000 629.350 499.560 ;
        RECT 630.040 499.500 630.360 499.560 ;
        RECT 628.750 497.860 629.350 498.000 ;
        RECT 628.750 497.040 628.890 497.860 ;
        RECT 628.430 496.840 628.890 497.040 ;
        RECT 628.430 496.780 628.750 496.840 ;
        RECT 628.430 17.580 628.750 17.640 ;
        RECT 2490.970 17.580 2491.290 17.640 ;
        RECT 628.430 17.440 2491.290 17.580 ;
        RECT 628.430 17.380 628.750 17.440 ;
        RECT 2490.970 17.380 2491.290 17.440 ;
      LAYER via ;
        RECT 630.070 499.500 630.330 499.760 ;
        RECT 628.460 496.780 628.720 497.040 ;
        RECT 628.460 17.380 628.720 17.640 ;
        RECT 2491.000 17.380 2491.260 17.640 ;
      LAYER met2 ;
        RECT 630.090 500.000 630.370 504.000 ;
        RECT 630.130 499.790 630.270 500.000 ;
        RECT 630.070 499.470 630.330 499.790 ;
        RECT 628.460 496.750 628.720 497.070 ;
        RECT 628.520 17.670 628.660 496.750 ;
        RECT 628.460 17.350 628.720 17.670 ;
        RECT 2491.000 17.350 2491.260 17.670 ;
        RECT 2491.060 2.400 2491.200 17.350 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.410 17.240 634.730 17.300 ;
        RECT 2508.910 17.240 2509.230 17.300 ;
        RECT 634.410 17.100 2509.230 17.240 ;
        RECT 634.410 17.040 634.730 17.100 ;
        RECT 2508.910 17.040 2509.230 17.100 ;
      LAYER via ;
        RECT 634.440 17.040 634.700 17.300 ;
        RECT 2508.940 17.040 2509.200 17.300 ;
      LAYER met2 ;
        RECT 631.470 500.000 631.750 504.000 ;
        RECT 631.510 499.475 631.650 500.000 ;
        RECT 631.440 499.105 631.720 499.475 ;
        RECT 634.430 497.235 634.710 497.605 ;
        RECT 634.500 17.330 634.640 497.235 ;
        RECT 634.440 17.010 634.700 17.330 ;
        RECT 2508.940 17.010 2509.200 17.330 ;
        RECT 2509.000 2.400 2509.140 17.010 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
      LAYER via2 ;
        RECT 631.440 499.150 631.720 499.430 ;
        RECT 634.430 497.280 634.710 497.560 ;
      LAYER met3 ;
        RECT 631.415 499.125 631.745 499.455 ;
        RECT 631.430 497.570 631.730 499.125 ;
        RECT 634.405 497.570 634.735 497.585 ;
        RECT 631.430 497.270 634.735 497.570 ;
        RECT 634.405 497.255 634.735 497.270 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.850 500.000 633.130 504.000 ;
        RECT 632.890 498.340 633.030 500.000 ;
        RECT 632.890 498.200 633.260 498.340 ;
        RECT 633.120 484.005 633.260 498.200 ;
        RECT 633.050 483.635 633.330 484.005 ;
        RECT 2526.870 16.475 2527.150 16.845 ;
        RECT 2526.940 2.400 2527.080 16.475 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
      LAYER via2 ;
        RECT 633.050 483.680 633.330 483.960 ;
        RECT 2526.870 16.520 2527.150 16.800 ;
      LAYER met3 ;
        RECT 633.025 483.970 633.355 483.985 ;
        RECT 634.150 483.970 634.530 483.980 ;
        RECT 633.025 483.670 634.530 483.970 ;
        RECT 633.025 483.655 633.355 483.670 ;
        RECT 634.150 483.660 634.530 483.670 ;
        RECT 634.150 16.810 634.530 16.820 ;
        RECT 2526.845 16.810 2527.175 16.825 ;
        RECT 634.150 16.510 2527.175 16.810 ;
        RECT 634.150 16.500 634.530 16.510 ;
        RECT 2526.845 16.495 2527.175 16.510 ;
      LAYER via3 ;
        RECT 634.180 483.660 634.500 483.980 ;
        RECT 634.180 16.500 634.500 16.820 ;
      LAYER met4 ;
        RECT 634.175 483.655 634.505 483.985 ;
        RECT 634.190 16.825 634.490 483.655 ;
        RECT 634.175 16.495 634.505 16.825 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 633.950 488.140 634.270 488.200 ;
        RECT 1928.390 488.140 1928.710 488.200 ;
        RECT 633.950 488.000 1928.710 488.140 ;
        RECT 633.950 487.940 634.270 488.000 ;
        RECT 1928.390 487.940 1928.710 488.000 ;
        RECT 1928.390 19.280 1928.710 19.340 ;
        RECT 2544.330 19.280 2544.650 19.340 ;
        RECT 1928.390 19.140 2544.650 19.280 ;
        RECT 1928.390 19.080 1928.710 19.140 ;
        RECT 2544.330 19.080 2544.650 19.140 ;
      LAYER via ;
        RECT 633.980 487.940 634.240 488.200 ;
        RECT 1928.420 487.940 1928.680 488.200 ;
        RECT 1928.420 19.080 1928.680 19.340 ;
        RECT 2544.360 19.080 2544.620 19.340 ;
      LAYER met2 ;
        RECT 634.230 500.000 634.510 504.000 ;
        RECT 634.270 499.645 634.410 500.000 ;
        RECT 634.200 499.275 634.480 499.645 ;
        RECT 633.970 498.595 634.250 498.965 ;
        RECT 634.040 488.230 634.180 498.595 ;
        RECT 633.980 487.910 634.240 488.230 ;
        RECT 1928.420 487.910 1928.680 488.230 ;
        RECT 1928.480 19.370 1928.620 487.910 ;
        RECT 1928.420 19.050 1928.680 19.370 ;
        RECT 2544.360 19.050 2544.620 19.370 ;
        RECT 2544.420 2.400 2544.560 19.050 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
      LAYER via2 ;
        RECT 634.200 499.320 634.480 499.600 ;
        RECT 633.970 498.640 634.250 498.920 ;
      LAYER met3 ;
        RECT 634.175 499.295 634.505 499.625 ;
        RECT 634.190 498.945 634.490 499.295 ;
        RECT 633.945 498.630 634.490 498.945 ;
        RECT 633.945 498.615 634.275 498.630 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 635.560 502.080 635.880 502.140 ;
        RECT 667.070 502.080 667.390 502.140 ;
        RECT 635.560 501.940 667.390 502.080 ;
        RECT 635.560 501.880 635.880 501.940 ;
        RECT 667.070 501.880 667.390 501.940 ;
        RECT 665.690 24.720 666.010 24.780 ;
        RECT 2562.270 24.720 2562.590 24.780 ;
        RECT 665.690 24.580 2562.590 24.720 ;
        RECT 665.690 24.520 666.010 24.580 ;
        RECT 2562.270 24.520 2562.590 24.580 ;
      LAYER via ;
        RECT 635.590 501.880 635.850 502.140 ;
        RECT 667.100 501.880 667.360 502.140 ;
        RECT 665.720 24.520 665.980 24.780 ;
        RECT 2562.300 24.520 2562.560 24.780 ;
      LAYER met2 ;
        RECT 635.610 502.170 635.890 504.000 ;
        RECT 635.590 501.850 635.890 502.170 ;
        RECT 667.100 501.850 667.360 502.170 ;
        RECT 635.610 500.000 635.890 501.850 ;
        RECT 667.160 489.330 667.300 501.850 ;
        RECT 665.320 489.190 667.300 489.330 ;
        RECT 665.320 448.570 665.460 489.190 ;
        RECT 665.320 448.430 665.920 448.570 ;
        RECT 665.780 24.810 665.920 448.430 ;
        RECT 665.720 24.490 665.980 24.810 ;
        RECT 2562.300 24.490 2562.560 24.810 ;
        RECT 2562.360 2.400 2562.500 24.490 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 800.930 489.500 801.250 489.560 ;
        RECT 548.710 489.360 801.250 489.500 ;
        RECT 517.110 489.160 517.430 489.220 ;
        RECT 548.710 489.160 548.850 489.360 ;
        RECT 800.930 489.300 801.250 489.360 ;
        RECT 517.110 489.020 548.850 489.160 ;
        RECT 517.110 488.960 517.430 489.020 ;
      LAYER via ;
        RECT 517.140 488.960 517.400 489.220 ;
        RECT 800.960 489.300 801.220 489.560 ;
      LAYER met2 ;
        RECT 498.990 500.000 499.270 504.000 ;
        RECT 499.030 499.645 499.170 500.000 ;
        RECT 498.960 499.275 499.240 499.645 ;
        RECT 517.130 489.075 517.410 489.445 ;
        RECT 800.960 489.270 801.220 489.590 ;
        RECT 517.140 488.930 517.400 489.075 ;
        RECT 801.020 82.870 801.160 489.270 ;
        RECT 801.020 82.730 806.680 82.870 ;
        RECT 806.540 2.400 806.680 82.730 ;
        RECT 806.330 -4.800 806.890 2.400 ;
      LAYER via2 ;
        RECT 498.960 499.320 499.240 499.600 ;
        RECT 517.130 489.120 517.410 489.400 ;
      LAYER met3 ;
        RECT 498.935 499.620 499.265 499.625 ;
        RECT 498.910 499.610 499.290 499.620 ;
        RECT 498.480 499.310 499.290 499.610 ;
        RECT 498.910 499.300 499.290 499.310 ;
        RECT 498.935 499.295 499.265 499.300 ;
        RECT 498.910 489.410 499.290 489.420 ;
        RECT 517.105 489.410 517.435 489.425 ;
        RECT 498.910 489.110 517.435 489.410 ;
        RECT 498.910 489.100 499.290 489.110 ;
        RECT 517.105 489.095 517.435 489.110 ;
      LAYER via3 ;
        RECT 498.940 499.300 499.260 499.620 ;
        RECT 498.940 489.100 499.260 489.420 ;
      LAYER met4 ;
        RECT 498.935 499.295 499.265 499.625 ;
        RECT 498.950 489.425 499.250 499.295 ;
        RECT 498.935 489.095 499.265 489.425 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 637.630 490.860 637.950 490.920 ;
        RECT 654.650 490.860 654.970 490.920 ;
        RECT 637.630 490.720 654.970 490.860 ;
        RECT 637.630 490.660 637.950 490.720 ;
        RECT 654.650 490.660 654.970 490.720 ;
        RECT 654.650 486.780 654.970 486.840 ;
        RECT 2573.770 486.780 2574.090 486.840 ;
        RECT 654.650 486.640 2574.090 486.780 ;
        RECT 654.650 486.580 654.970 486.640 ;
        RECT 2573.770 486.580 2574.090 486.640 ;
        RECT 2573.770 17.580 2574.090 17.640 ;
        RECT 2577.910 17.580 2578.230 17.640 ;
        RECT 2573.770 17.440 2578.230 17.580 ;
        RECT 2573.770 17.380 2574.090 17.440 ;
        RECT 2577.910 17.380 2578.230 17.440 ;
      LAYER via ;
        RECT 637.660 490.660 637.920 490.920 ;
        RECT 654.680 490.660 654.940 490.920 ;
        RECT 654.680 486.580 654.940 486.840 ;
        RECT 2573.800 486.580 2574.060 486.840 ;
        RECT 2573.800 17.380 2574.060 17.640 ;
        RECT 2577.940 17.380 2578.200 17.640 ;
      LAYER met2 ;
        RECT 636.990 500.000 637.270 504.000 ;
        RECT 637.030 499.645 637.170 500.000 ;
        RECT 636.960 499.275 637.240 499.645 ;
        RECT 637.650 498.595 637.930 498.965 ;
        RECT 637.720 490.950 637.860 498.595 ;
        RECT 637.660 490.630 637.920 490.950 ;
        RECT 654.680 490.630 654.940 490.950 ;
        RECT 654.740 486.870 654.880 490.630 ;
        RECT 654.680 486.550 654.940 486.870 ;
        RECT 2573.800 486.550 2574.060 486.870 ;
        RECT 2573.860 17.670 2574.000 486.550 ;
        RECT 2573.800 17.350 2574.060 17.670 ;
        RECT 2577.940 17.350 2578.200 17.670 ;
        RECT 2578.000 1.770 2578.140 17.350 ;
        RECT 2579.630 1.770 2580.190 2.400 ;
        RECT 2578.000 1.630 2580.190 1.770 ;
        RECT 2579.630 -4.800 2580.190 1.630 ;
      LAYER via2 ;
        RECT 636.960 499.320 637.240 499.600 ;
        RECT 637.650 498.640 637.930 498.920 ;
      LAYER met3 ;
        RECT 636.935 499.295 637.265 499.625 ;
        RECT 636.950 498.930 637.250 499.295 ;
        RECT 637.625 498.930 637.955 498.945 ;
        RECT 636.950 498.630 637.955 498.930 ;
        RECT 637.625 498.615 637.955 498.630 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.370 500.000 638.650 504.000 ;
        RECT 669.390 500.635 669.670 501.005 ;
        RECT 638.410 499.815 638.550 500.000 ;
        RECT 638.340 499.445 638.620 499.815 ;
        RECT 669.460 486.045 669.600 500.635 ;
        RECT 669.390 485.675 669.670 486.045 ;
        RECT 2594.490 485.675 2594.770 486.045 ;
        RECT 2594.560 82.870 2594.700 485.675 ;
        RECT 2594.560 82.730 2597.920 82.870 ;
        RECT 2597.780 2.400 2597.920 82.730 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
      LAYER via2 ;
        RECT 669.390 500.680 669.670 500.960 ;
        RECT 638.340 499.490 638.620 499.770 ;
        RECT 669.390 485.720 669.670 486.000 ;
        RECT 2594.490 485.720 2594.770 486.000 ;
      LAYER met3 ;
        RECT 669.365 500.970 669.695 500.985 ;
        RECT 638.330 500.670 669.695 500.970 ;
        RECT 638.330 499.795 638.630 500.670 ;
        RECT 669.365 500.655 669.695 500.670 ;
        RECT 638.315 499.465 638.645 499.795 ;
        RECT 669.365 486.010 669.695 486.025 ;
        RECT 2594.465 486.010 2594.795 486.025 ;
        RECT 669.365 485.710 2594.795 486.010 ;
        RECT 669.365 485.695 669.695 485.710 ;
        RECT 2594.465 485.695 2594.795 485.710 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 639.700 499.500 640.020 499.760 ;
        RECT 639.790 498.060 639.930 499.500 ;
        RECT 639.790 497.860 640.250 498.060 ;
        RECT 639.930 497.800 640.250 497.860 ;
        RECT 634.870 471.140 635.190 471.200 ;
        RECT 639.470 471.140 639.790 471.200 ;
        RECT 634.870 471.000 639.790 471.140 ;
        RECT 634.870 470.940 635.190 471.000 ;
        RECT 639.470 470.940 639.790 471.000 ;
        RECT 634.870 24.380 635.190 24.440 ;
        RECT 2615.170 24.380 2615.490 24.440 ;
        RECT 634.870 24.240 2615.490 24.380 ;
        RECT 634.870 24.180 635.190 24.240 ;
        RECT 2615.170 24.180 2615.490 24.240 ;
      LAYER via ;
        RECT 639.730 499.500 639.990 499.760 ;
        RECT 639.960 497.800 640.220 498.060 ;
        RECT 634.900 470.940 635.160 471.200 ;
        RECT 639.500 470.940 639.760 471.200 ;
        RECT 634.900 24.180 635.160 24.440 ;
        RECT 2615.200 24.180 2615.460 24.440 ;
      LAYER met2 ;
        RECT 639.750 500.000 640.030 504.000 ;
        RECT 639.790 499.790 639.930 500.000 ;
        RECT 639.730 499.470 639.990 499.790 ;
        RECT 639.960 497.770 640.220 498.090 ;
        RECT 640.020 489.970 640.160 497.770 ;
        RECT 639.560 489.830 640.160 489.970 ;
        RECT 639.560 471.230 639.700 489.830 ;
        RECT 634.900 470.910 635.160 471.230 ;
        RECT 639.500 470.910 639.760 471.230 ;
        RECT 634.960 24.470 635.100 470.910 ;
        RECT 634.900 24.150 635.160 24.470 ;
        RECT 2615.200 24.150 2615.460 24.470 ;
        RECT 2615.260 2.400 2615.400 24.150 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 641.080 499.160 641.400 499.420 ;
        RECT 641.170 498.400 641.310 499.160 ;
        RECT 640.850 498.200 641.310 498.400 ;
        RECT 640.850 498.140 641.170 498.200 ;
      LAYER via ;
        RECT 641.110 499.160 641.370 499.420 ;
        RECT 640.880 498.140 641.140 498.400 ;
      LAYER met2 ;
        RECT 641.130 500.000 641.410 504.000 ;
        RECT 641.170 499.450 641.310 500.000 ;
        RECT 641.110 499.130 641.370 499.450 ;
        RECT 640.880 498.110 641.140 498.430 ;
        RECT 640.940 487.405 641.080 498.110 ;
        RECT 640.870 487.035 641.150 487.405 ;
        RECT 2633.130 25.995 2633.410 26.365 ;
        RECT 2633.200 2.400 2633.340 25.995 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
      LAYER via2 ;
        RECT 640.870 487.080 641.150 487.360 ;
        RECT 2633.130 26.040 2633.410 26.320 ;
      LAYER met3 ;
        RECT 637.830 487.370 638.210 487.380 ;
        RECT 640.845 487.370 641.175 487.385 ;
        RECT 637.830 487.070 641.175 487.370 ;
        RECT 637.830 487.060 638.210 487.070 ;
        RECT 640.845 487.055 641.175 487.070 ;
        RECT 637.830 26.330 638.210 26.340 ;
        RECT 2633.105 26.330 2633.435 26.345 ;
        RECT 637.830 26.030 2633.435 26.330 ;
        RECT 637.830 26.020 638.210 26.030 ;
        RECT 2633.105 26.015 2633.435 26.030 ;
      LAYER via3 ;
        RECT 637.860 487.060 638.180 487.380 ;
        RECT 637.860 26.020 638.180 26.340 ;
      LAYER met4 ;
        RECT 637.855 487.055 638.185 487.385 ;
        RECT 637.870 26.345 638.170 487.055 ;
        RECT 637.855 26.015 638.185 26.345 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 642.460 499.160 642.780 499.420 ;
        RECT 642.550 496.980 642.690 499.160 ;
        RECT 662.930 496.980 663.250 497.040 ;
        RECT 642.550 496.840 663.250 496.980 ;
        RECT 662.930 496.780 663.250 496.840 ;
        RECT 662.930 493.240 663.250 493.300 ;
        RECT 2649.670 493.240 2649.990 493.300 ;
        RECT 662.930 493.100 2649.990 493.240 ;
        RECT 662.930 493.040 663.250 493.100 ;
        RECT 2649.670 493.040 2649.990 493.100 ;
      LAYER via ;
        RECT 642.490 499.160 642.750 499.420 ;
        RECT 662.960 496.780 663.220 497.040 ;
        RECT 662.960 493.040 663.220 493.300 ;
        RECT 2649.700 493.040 2649.960 493.300 ;
      LAYER met2 ;
        RECT 642.510 500.000 642.790 504.000 ;
        RECT 642.550 499.450 642.690 500.000 ;
        RECT 642.490 499.130 642.750 499.450 ;
        RECT 662.960 496.750 663.220 497.070 ;
        RECT 663.020 493.330 663.160 496.750 ;
        RECT 662.960 493.010 663.220 493.330 ;
        RECT 2649.700 493.010 2649.960 493.330 ;
        RECT 2649.760 1.770 2649.900 493.010 ;
        RECT 2650.470 1.770 2651.030 2.400 ;
        RECT 2649.760 1.630 2651.030 1.770 ;
        RECT 2650.470 -4.800 2651.030 1.630 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 643.840 499.160 644.160 499.420 ;
        RECT 643.930 498.740 644.070 499.160 ;
        RECT 643.930 498.540 644.390 498.740 ;
        RECT 644.070 498.480 644.390 498.540 ;
        RECT 642.690 489.840 643.010 489.900 ;
        RECT 643.610 489.840 643.930 489.900 ;
        RECT 642.690 489.700 643.930 489.840 ;
        RECT 642.690 489.640 643.010 489.700 ;
        RECT 643.610 489.640 643.930 489.700 ;
        RECT 642.690 32.540 643.010 32.600 ;
        RECT 2668.530 32.540 2668.850 32.600 ;
        RECT 642.690 32.400 2668.850 32.540 ;
        RECT 642.690 32.340 643.010 32.400 ;
        RECT 2668.530 32.340 2668.850 32.400 ;
      LAYER via ;
        RECT 643.870 499.160 644.130 499.420 ;
        RECT 644.100 498.480 644.360 498.740 ;
        RECT 642.720 489.640 642.980 489.900 ;
        RECT 643.640 489.640 643.900 489.900 ;
        RECT 642.720 32.340 642.980 32.600 ;
        RECT 2668.560 32.340 2668.820 32.600 ;
      LAYER met2 ;
        RECT 643.890 500.000 644.170 504.000 ;
        RECT 643.930 499.450 644.070 500.000 ;
        RECT 643.870 499.130 644.130 499.450 ;
        RECT 644.100 498.450 644.360 498.770 ;
        RECT 644.160 498.170 644.300 498.450 ;
        RECT 643.700 498.030 644.300 498.170 ;
        RECT 643.700 489.930 643.840 498.030 ;
        RECT 642.720 489.610 642.980 489.930 ;
        RECT 643.640 489.610 643.900 489.930 ;
        RECT 642.780 32.630 642.920 489.610 ;
        RECT 642.720 32.310 642.980 32.630 ;
        RECT 2668.560 32.310 2668.820 32.630 ;
        RECT 2668.620 2.400 2668.760 32.310 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 642.230 487.460 642.550 487.520 ;
        RECT 645.450 487.460 645.770 487.520 ;
        RECT 642.230 487.320 645.770 487.460 ;
        RECT 642.230 487.260 642.550 487.320 ;
        RECT 645.450 487.260 645.770 487.320 ;
        RECT 642.230 31.860 642.550 31.920 ;
        RECT 2686.010 31.860 2686.330 31.920 ;
        RECT 642.230 31.720 2686.330 31.860 ;
        RECT 642.230 31.660 642.550 31.720 ;
        RECT 2686.010 31.660 2686.330 31.720 ;
      LAYER via ;
        RECT 642.260 487.260 642.520 487.520 ;
        RECT 645.480 487.260 645.740 487.520 ;
        RECT 642.260 31.660 642.520 31.920 ;
        RECT 2686.040 31.660 2686.300 31.920 ;
      LAYER met2 ;
        RECT 645.270 500.000 645.550 504.000 ;
        RECT 645.310 498.000 645.450 500.000 ;
        RECT 645.310 497.860 645.680 498.000 ;
        RECT 645.540 487.550 645.680 497.860 ;
        RECT 642.260 487.230 642.520 487.550 ;
        RECT 645.480 487.230 645.740 487.550 ;
        RECT 642.320 31.950 642.460 487.230 ;
        RECT 642.260 31.630 642.520 31.950 ;
        RECT 2686.040 31.630 2686.300 31.950 ;
        RECT 2686.100 2.400 2686.240 31.630 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 646.600 499.360 646.920 499.420 ;
        RECT 646.230 499.220 646.920 499.360 ;
        RECT 646.230 498.400 646.370 499.220 ;
        RECT 646.600 499.160 646.920 499.220 ;
        RECT 646.230 498.200 646.690 498.400 ;
        RECT 646.370 498.140 646.690 498.200 ;
        RECT 643.610 31.520 643.930 31.580 ;
        RECT 2703.950 31.520 2704.270 31.580 ;
        RECT 643.610 31.380 2704.270 31.520 ;
        RECT 643.610 31.320 643.930 31.380 ;
        RECT 2703.950 31.320 2704.270 31.380 ;
      LAYER via ;
        RECT 646.630 499.160 646.890 499.420 ;
        RECT 646.400 498.140 646.660 498.400 ;
        RECT 643.640 31.320 643.900 31.580 ;
        RECT 2703.980 31.320 2704.240 31.580 ;
      LAYER met2 ;
        RECT 646.650 500.000 646.930 504.000 ;
        RECT 646.690 499.450 646.830 500.000 ;
        RECT 646.630 499.130 646.890 499.450 ;
        RECT 646.400 498.285 646.660 498.430 ;
        RECT 646.390 497.915 646.670 498.285 ;
        RECT 644.090 497.235 644.370 497.605 ;
        RECT 644.160 473.010 644.300 497.235 ;
        RECT 643.700 472.870 644.300 473.010 ;
        RECT 643.700 31.610 643.840 472.870 ;
        RECT 643.640 31.290 643.900 31.610 ;
        RECT 2703.980 31.290 2704.240 31.610 ;
        RECT 2704.040 2.400 2704.180 31.290 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
      LAYER via2 ;
        RECT 646.390 497.960 646.670 498.240 ;
        RECT 644.090 497.280 644.370 497.560 ;
      LAYER met3 ;
        RECT 646.365 498.250 646.695 498.265 ;
        RECT 646.150 497.935 646.695 498.250 ;
        RECT 644.065 497.570 644.395 497.585 ;
        RECT 646.150 497.570 646.450 497.935 ;
        RECT 644.065 497.270 646.450 497.570 ;
        RECT 644.065 497.255 644.395 497.270 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.030 500.000 648.310 504.000 ;
        RECT 648.070 498.965 648.210 500.000 ;
        RECT 648.000 498.595 648.280 498.965 ;
        RECT 2721.910 30.755 2722.190 31.125 ;
        RECT 2721.980 2.400 2722.120 30.755 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
      LAYER via2 ;
        RECT 648.000 498.640 648.280 498.920 ;
        RECT 2721.910 30.800 2722.190 31.080 ;
      LAYER met3 ;
        RECT 647.975 498.940 648.305 498.945 ;
        RECT 647.950 498.930 648.330 498.940 ;
        RECT 647.520 498.630 648.330 498.930 ;
        RECT 647.950 498.620 648.330 498.630 ;
        RECT 647.975 498.615 648.305 498.620 ;
        RECT 647.950 31.090 648.330 31.100 ;
        RECT 2721.885 31.090 2722.215 31.105 ;
        RECT 647.950 30.790 2722.215 31.090 ;
        RECT 647.950 30.780 648.330 30.790 ;
        RECT 2721.885 30.775 2722.215 30.790 ;
      LAYER via3 ;
        RECT 647.980 498.620 648.300 498.940 ;
        RECT 647.980 30.780 648.300 31.100 ;
      LAYER met4 ;
        RECT 647.975 498.615 648.305 498.945 ;
        RECT 647.990 31.105 648.290 498.615 ;
        RECT 647.975 30.775 648.305 31.105 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 649.360 499.700 649.680 499.760 ;
        RECT 648.300 499.560 649.680 499.700 ;
        RECT 648.300 498.060 648.440 499.560 ;
        RECT 649.360 499.500 649.680 499.560 ;
        RECT 648.210 497.800 648.530 498.060 ;
      LAYER via ;
        RECT 649.390 499.500 649.650 499.760 ;
        RECT 648.240 497.800 648.500 498.060 ;
      LAYER met2 ;
        RECT 649.410 500.000 649.690 504.000 ;
        RECT 649.450 499.790 649.590 500.000 ;
        RECT 649.390 499.470 649.650 499.790 ;
        RECT 648.240 497.770 648.500 498.090 ;
        RECT 648.300 497.605 648.440 497.770 ;
        RECT 648.230 497.235 648.510 497.605 ;
        RECT 2739.390 493.155 2739.670 493.525 ;
        RECT 2739.460 2.400 2739.600 493.155 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
      LAYER via2 ;
        RECT 648.230 497.280 648.510 497.560 ;
        RECT 2739.390 493.200 2739.670 493.480 ;
      LAYER met3 ;
        RECT 648.205 497.570 648.535 497.585 ;
        RECT 648.870 497.570 649.250 497.580 ;
        RECT 648.205 497.270 649.250 497.570 ;
        RECT 648.205 497.255 648.535 497.270 ;
        RECT 648.870 497.260 649.250 497.270 ;
        RECT 648.870 493.490 649.250 493.500 ;
        RECT 2739.365 493.490 2739.695 493.505 ;
        RECT 648.870 493.190 2739.695 493.490 ;
        RECT 648.870 493.180 649.250 493.190 ;
        RECT 2739.365 493.175 2739.695 493.190 ;
      LAYER via3 ;
        RECT 648.900 497.260 649.220 497.580 ;
        RECT 648.900 493.180 649.220 493.500 ;
      LAYER met4 ;
        RECT 648.895 497.255 649.225 497.585 ;
        RECT 648.910 493.505 649.210 497.255 ;
        RECT 648.895 493.175 649.225 493.505 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 500.320 499.160 500.640 499.420 ;
        RECT 500.410 498.000 500.550 499.160 ;
        RECT 497.880 497.860 500.550 498.000 ;
        RECT 497.880 497.720 498.020 497.860 ;
        RECT 497.790 497.460 498.110 497.720 ;
        RECT 497.790 41.380 498.110 41.440 ;
        RECT 824.390 41.380 824.710 41.440 ;
        RECT 497.790 41.240 824.710 41.380 ;
        RECT 497.790 41.180 498.110 41.240 ;
        RECT 824.390 41.180 824.710 41.240 ;
      LAYER via ;
        RECT 500.350 499.160 500.610 499.420 ;
        RECT 497.820 497.460 498.080 497.720 ;
        RECT 497.820 41.180 498.080 41.440 ;
        RECT 824.420 41.180 824.680 41.440 ;
      LAYER met2 ;
        RECT 500.370 500.000 500.650 504.000 ;
        RECT 500.410 499.450 500.550 500.000 ;
        RECT 500.350 499.130 500.610 499.450 ;
        RECT 497.820 497.430 498.080 497.750 ;
        RECT 497.880 41.470 498.020 497.430 ;
        RECT 497.820 41.150 498.080 41.470 ;
        RECT 824.420 41.150 824.680 41.470 ;
        RECT 824.480 2.400 824.620 41.150 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 650.740 499.500 651.060 499.760 ;
        RECT 650.830 498.680 650.970 499.500 ;
        RECT 650.370 498.540 650.970 498.680 ;
        RECT 650.370 498.000 650.510 498.540 ;
        RECT 650.970 498.000 651.290 498.060 ;
        RECT 650.370 497.860 651.290 498.000 ;
        RECT 650.970 497.800 651.290 497.860 ;
        RECT 649.590 472.840 649.910 472.900 ;
        RECT 650.970 472.840 651.290 472.900 ;
        RECT 649.590 472.700 651.290 472.840 ;
        RECT 649.590 472.640 649.910 472.700 ;
        RECT 650.970 472.640 651.290 472.700 ;
        RECT 649.590 39.680 649.910 39.740 ;
        RECT 2757.310 39.680 2757.630 39.740 ;
        RECT 649.590 39.540 2757.630 39.680 ;
        RECT 649.590 39.480 649.910 39.540 ;
        RECT 2757.310 39.480 2757.630 39.540 ;
      LAYER via ;
        RECT 650.770 499.500 651.030 499.760 ;
        RECT 651.000 497.800 651.260 498.060 ;
        RECT 649.620 472.640 649.880 472.900 ;
        RECT 651.000 472.640 651.260 472.900 ;
        RECT 649.620 39.480 649.880 39.740 ;
        RECT 2757.340 39.480 2757.600 39.740 ;
      LAYER met2 ;
        RECT 650.790 500.000 651.070 504.000 ;
        RECT 650.830 499.790 650.970 500.000 ;
        RECT 650.770 499.470 651.030 499.790 ;
        RECT 651.000 497.770 651.260 498.090 ;
        RECT 651.060 472.930 651.200 497.770 ;
        RECT 649.620 472.610 649.880 472.930 ;
        RECT 651.000 472.610 651.260 472.930 ;
        RECT 649.680 39.770 649.820 472.610 ;
        RECT 649.620 39.450 649.880 39.770 ;
        RECT 2757.340 39.450 2757.600 39.770 ;
        RECT 2757.400 2.400 2757.540 39.450 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 652.120 499.500 652.440 499.760 ;
        RECT 652.210 499.360 652.350 499.500 ;
        RECT 652.210 499.220 652.580 499.360 ;
        RECT 650.050 497.320 650.370 497.380 ;
        RECT 652.440 497.320 652.580 499.220 ;
        RECT 650.050 497.180 652.580 497.320 ;
        RECT 650.050 497.120 650.370 497.180 ;
        RECT 650.050 474.880 650.370 474.940 ;
        RECT 648.760 474.740 650.370 474.880 ;
        RECT 648.760 473.240 648.900 474.740 ;
        RECT 650.050 474.680 650.370 474.740 ;
        RECT 648.670 472.980 648.990 473.240 ;
        RECT 648.670 24.040 648.990 24.100 ;
        RECT 2774.790 24.040 2775.110 24.100 ;
        RECT 648.670 23.900 2775.110 24.040 ;
        RECT 648.670 23.840 648.990 23.900 ;
        RECT 2774.790 23.840 2775.110 23.900 ;
      LAYER via ;
        RECT 652.150 499.500 652.410 499.760 ;
        RECT 650.080 497.120 650.340 497.380 ;
        RECT 650.080 474.680 650.340 474.940 ;
        RECT 648.700 472.980 648.960 473.240 ;
        RECT 648.700 23.840 648.960 24.100 ;
        RECT 2774.820 23.840 2775.080 24.100 ;
      LAYER met2 ;
        RECT 652.170 500.000 652.450 504.000 ;
        RECT 652.210 499.790 652.350 500.000 ;
        RECT 652.150 499.470 652.410 499.790 ;
        RECT 650.080 497.090 650.340 497.410 ;
        RECT 650.140 474.970 650.280 497.090 ;
        RECT 650.080 474.650 650.340 474.970 ;
        RECT 648.700 472.950 648.960 473.270 ;
        RECT 648.760 24.130 648.900 472.950 ;
        RECT 648.700 23.810 648.960 24.130 ;
        RECT 2774.820 23.810 2775.080 24.130 ;
        RECT 2774.880 2.400 2775.020 23.810 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.550 500.000 653.830 504.000 ;
        RECT 653.590 499.815 653.730 500.000 ;
        RECT 653.520 499.445 653.800 499.815 ;
        RECT 2792.750 25.315 2793.030 25.685 ;
        RECT 2792.820 2.400 2792.960 25.315 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
      LAYER via2 ;
        RECT 653.520 499.490 653.800 499.770 ;
        RECT 2792.750 25.360 2793.030 25.640 ;
      LAYER met3 ;
        RECT 653.495 499.465 653.825 499.795 ;
        RECT 653.510 498.940 653.810 499.465 ;
        RECT 653.470 498.620 653.850 498.940 ;
        RECT 653.470 25.650 653.850 25.660 ;
        RECT 2792.725 25.650 2793.055 25.665 ;
        RECT 653.470 25.350 2793.055 25.650 ;
        RECT 653.470 25.340 653.850 25.350 ;
        RECT 2792.725 25.335 2793.055 25.350 ;
      LAYER via3 ;
        RECT 653.500 498.620 653.820 498.940 ;
        RECT 653.500 25.340 653.820 25.660 ;
      LAYER met4 ;
        RECT 653.495 498.615 653.825 498.945 ;
        RECT 653.510 25.665 653.810 498.615 ;
        RECT 653.495 25.335 653.825 25.665 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 654.880 499.160 655.200 499.420 ;
        RECT 654.970 498.400 655.110 499.160 ;
        RECT 654.970 498.200 655.430 498.400 ;
        RECT 655.110 498.140 655.430 498.200 ;
      LAYER via ;
        RECT 654.910 499.160 655.170 499.420 ;
        RECT 655.140 498.140 655.400 498.400 ;
      LAYER met2 ;
        RECT 654.930 500.000 655.210 504.000 ;
        RECT 654.970 499.450 655.110 500.000 ;
        RECT 654.910 499.130 655.170 499.450 ;
        RECT 655.140 498.110 655.400 498.430 ;
        RECT 655.200 494.885 655.340 498.110 ;
        RECT 655.130 494.515 655.410 494.885 ;
        RECT 2810.230 24.635 2810.510 25.005 ;
        RECT 2810.300 2.400 2810.440 24.635 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
      LAYER via2 ;
        RECT 655.130 494.560 655.410 494.840 ;
        RECT 2810.230 24.680 2810.510 24.960 ;
      LAYER met3 ;
        RECT 654.390 494.850 654.770 494.860 ;
        RECT 655.105 494.850 655.435 494.865 ;
        RECT 654.390 494.550 655.435 494.850 ;
        RECT 654.390 494.540 654.770 494.550 ;
        RECT 655.105 494.535 655.435 494.550 ;
        RECT 654.390 24.970 654.770 24.980 ;
        RECT 2810.205 24.970 2810.535 24.985 ;
        RECT 654.390 24.670 2810.535 24.970 ;
        RECT 654.390 24.660 654.770 24.670 ;
        RECT 2810.205 24.655 2810.535 24.670 ;
      LAYER via3 ;
        RECT 654.420 494.540 654.740 494.860 ;
        RECT 654.420 24.660 654.740 24.980 ;
      LAYER met4 ;
        RECT 654.415 494.535 654.745 494.865 ;
        RECT 654.430 24.985 654.730 494.535 ;
        RECT 654.415 24.655 654.745 24.985 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.260 499.500 656.580 499.760 ;
        RECT 656.350 498.740 656.490 499.500 ;
        RECT 656.350 498.540 656.810 498.740 ;
        RECT 656.490 498.480 656.810 498.540 ;
        RECT 656.950 39.340 657.270 39.400 ;
        RECT 2828.150 39.340 2828.470 39.400 ;
        RECT 656.950 39.200 2828.470 39.340 ;
        RECT 656.950 39.140 657.270 39.200 ;
        RECT 2828.150 39.140 2828.470 39.200 ;
      LAYER via ;
        RECT 656.290 499.500 656.550 499.760 ;
        RECT 656.520 498.480 656.780 498.740 ;
        RECT 656.980 39.140 657.240 39.400 ;
        RECT 2828.180 39.140 2828.440 39.400 ;
      LAYER met2 ;
        RECT 656.310 500.000 656.590 504.000 ;
        RECT 656.350 499.790 656.490 500.000 ;
        RECT 656.290 499.470 656.550 499.790 ;
        RECT 656.520 498.450 656.780 498.770 ;
        RECT 656.580 489.330 656.720 498.450 ;
        RECT 656.580 489.190 657.180 489.330 ;
        RECT 657.040 39.430 657.180 489.190 ;
        RECT 656.980 39.110 657.240 39.430 ;
        RECT 2828.180 39.110 2828.440 39.430 ;
        RECT 2828.240 2.400 2828.380 39.110 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 657.640 499.160 657.960 499.420 ;
        RECT 657.730 498.060 657.870 499.160 ;
        RECT 657.730 497.860 658.190 498.060 ;
        RECT 657.870 497.800 658.190 497.860 ;
        RECT 657.870 39.000 658.190 39.060 ;
        RECT 2845.630 39.000 2845.950 39.060 ;
        RECT 657.870 38.860 2845.950 39.000 ;
        RECT 657.870 38.800 658.190 38.860 ;
        RECT 2845.630 38.800 2845.950 38.860 ;
      LAYER via ;
        RECT 657.670 499.160 657.930 499.420 ;
        RECT 657.900 497.800 658.160 498.060 ;
        RECT 657.900 38.800 658.160 39.060 ;
        RECT 2845.660 38.800 2845.920 39.060 ;
      LAYER met2 ;
        RECT 657.690 500.000 657.970 504.000 ;
        RECT 657.730 499.450 657.870 500.000 ;
        RECT 657.670 499.130 657.930 499.450 ;
        RECT 657.900 497.770 658.160 498.090 ;
        RECT 657.960 39.090 658.100 497.770 ;
        RECT 657.900 38.770 658.160 39.090 ;
        RECT 2845.660 38.770 2845.920 39.090 ;
        RECT 2845.720 2.400 2845.860 38.770 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.030 471.820 656.350 471.880 ;
        RECT 661.550 471.820 661.870 471.880 ;
        RECT 656.030 471.680 661.870 471.820 ;
        RECT 656.030 471.620 656.350 471.680 ;
        RECT 661.550 471.620 661.870 471.680 ;
        RECT 656.030 37.980 656.350 38.040 ;
        RECT 2863.570 37.980 2863.890 38.040 ;
        RECT 656.030 37.840 2863.890 37.980 ;
        RECT 656.030 37.780 656.350 37.840 ;
        RECT 2863.570 37.780 2863.890 37.840 ;
      LAYER via ;
        RECT 656.060 471.620 656.320 471.880 ;
        RECT 661.580 471.620 661.840 471.880 ;
        RECT 656.060 37.780 656.320 38.040 ;
        RECT 2863.600 37.780 2863.860 38.040 ;
      LAYER met2 ;
        RECT 659.070 500.000 659.350 504.000 ;
        RECT 659.110 499.645 659.250 500.000 ;
        RECT 659.040 499.275 659.320 499.645 ;
        RECT 661.110 497.915 661.390 498.285 ;
        RECT 661.180 476.170 661.320 497.915 ;
        RECT 661.180 476.030 661.780 476.170 ;
        RECT 661.640 471.910 661.780 476.030 ;
        RECT 656.060 471.590 656.320 471.910 ;
        RECT 661.580 471.590 661.840 471.910 ;
        RECT 656.120 38.070 656.260 471.590 ;
        RECT 656.060 37.750 656.320 38.070 ;
        RECT 2863.600 37.750 2863.860 38.070 ;
        RECT 2863.660 2.400 2863.800 37.750 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
      LAYER via2 ;
        RECT 659.040 499.320 659.320 499.600 ;
        RECT 661.110 497.960 661.390 498.240 ;
      LAYER met3 ;
        RECT 659.015 499.295 659.345 499.625 ;
        RECT 659.030 498.250 659.330 499.295 ;
        RECT 661.085 498.250 661.415 498.265 ;
        RECT 659.030 497.950 661.415 498.250 ;
        RECT 661.085 497.935 661.415 497.950 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 660.400 499.160 660.720 499.420 ;
        RECT 660.490 498.680 660.630 499.160 ;
        RECT 660.260 498.540 660.630 498.680 ;
        RECT 660.260 498.060 660.400 498.540 ;
        RECT 660.170 497.800 660.490 498.060 ;
      LAYER via ;
        RECT 660.430 499.160 660.690 499.420 ;
        RECT 660.200 497.800 660.460 498.060 ;
      LAYER met2 ;
        RECT 660.450 500.000 660.730 504.000 ;
        RECT 660.490 499.450 660.630 500.000 ;
        RECT 660.430 499.130 660.690 499.450 ;
        RECT 660.200 497.770 660.460 498.090 ;
        RECT 660.260 490.805 660.400 497.770 ;
        RECT 660.190 490.435 660.470 490.805 ;
        RECT 2881.530 23.955 2881.810 24.325 ;
        RECT 2881.600 2.400 2881.740 23.955 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
      LAYER via2 ;
        RECT 660.190 490.480 660.470 490.760 ;
        RECT 2881.530 24.000 2881.810 24.280 ;
      LAYER met3 ;
        RECT 660.165 490.780 660.495 490.785 ;
        RECT 659.910 490.770 660.495 490.780 ;
        RECT 659.710 490.470 660.495 490.770 ;
        RECT 659.910 490.460 660.495 490.470 ;
        RECT 660.165 490.455 660.495 490.460 ;
        RECT 659.910 24.290 660.290 24.300 ;
        RECT 2881.505 24.290 2881.835 24.305 ;
        RECT 659.910 23.990 2881.835 24.290 ;
        RECT 659.910 23.980 660.290 23.990 ;
        RECT 2881.505 23.975 2881.835 23.990 ;
      LAYER via3 ;
        RECT 659.940 490.460 660.260 490.780 ;
        RECT 659.940 23.980 660.260 24.300 ;
      LAYER met4 ;
        RECT 659.935 490.455 660.265 490.785 ;
        RECT 659.950 24.305 660.250 490.455 ;
        RECT 659.935 23.975 660.265 24.305 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.750 500.000 502.030 504.000 ;
        RECT 501.790 499.645 501.930 500.000 ;
        RECT 501.720 499.275 502.000 499.645 ;
        RECT 842.350 45.035 842.630 45.405 ;
        RECT 842.420 17.410 842.560 45.035 ;
        RECT 841.960 17.270 842.560 17.410 ;
        RECT 841.960 2.400 842.100 17.270 ;
        RECT 841.750 -4.800 842.310 2.400 ;
      LAYER via2 ;
        RECT 501.720 499.320 502.000 499.600 ;
        RECT 842.350 45.080 842.630 45.360 ;
      LAYER met3 ;
        RECT 501.695 499.610 502.025 499.625 ;
        RECT 501.695 499.295 502.240 499.610 ;
        RECT 501.940 498.930 502.240 499.295 ;
        RECT 502.590 498.930 502.970 498.940 ;
        RECT 501.940 498.630 502.970 498.930 ;
        RECT 502.590 498.620 502.970 498.630 ;
        RECT 502.590 45.370 502.970 45.380 ;
        RECT 842.325 45.370 842.655 45.385 ;
        RECT 502.590 45.070 842.655 45.370 ;
        RECT 502.590 45.060 502.970 45.070 ;
        RECT 842.325 45.055 842.655 45.070 ;
      LAYER via3 ;
        RECT 502.620 498.620 502.940 498.940 ;
        RECT 502.620 45.060 502.940 45.380 ;
      LAYER met4 ;
        RECT 502.615 498.615 502.945 498.945 ;
        RECT 502.630 45.385 502.930 498.615 ;
        RECT 502.615 45.055 502.945 45.385 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.130 500.000 503.410 504.000 ;
        RECT 503.170 499.645 503.310 500.000 ;
        RECT 503.100 499.275 503.380 499.645 ;
        RECT 859.830 44.355 860.110 44.725 ;
        RECT 859.900 2.400 860.040 44.355 ;
        RECT 859.690 -4.800 860.250 2.400 ;
      LAYER via2 ;
        RECT 503.100 499.320 503.380 499.600 ;
        RECT 859.830 44.400 860.110 44.680 ;
      LAYER met3 ;
        RECT 501.670 500.290 502.050 500.300 ;
        RECT 501.670 499.990 503.160 500.290 ;
        RECT 501.670 499.980 502.050 499.990 ;
        RECT 502.860 499.625 503.160 499.990 ;
        RECT 502.860 499.310 503.405 499.625 ;
        RECT 503.075 499.295 503.405 499.310 ;
        RECT 501.670 44.690 502.050 44.700 ;
        RECT 859.805 44.690 860.135 44.705 ;
        RECT 501.670 44.390 860.135 44.690 ;
        RECT 501.670 44.380 502.050 44.390 ;
        RECT 859.805 44.375 860.135 44.390 ;
      LAYER via3 ;
        RECT 501.700 499.980 502.020 500.300 ;
        RECT 501.700 44.380 502.020 44.700 ;
      LAYER met4 ;
        RECT 501.695 499.975 502.025 500.305 ;
        RECT 501.710 44.705 502.010 499.975 ;
        RECT 501.695 44.375 502.025 44.705 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 570.470 490.520 570.790 490.580 ;
        RECT 531.230 490.380 570.790 490.520 ;
        RECT 504.690 489.840 505.010 489.900 ;
        RECT 531.230 489.840 531.370 490.380 ;
        RECT 570.470 490.320 570.790 490.380 ;
        RECT 504.690 489.700 531.370 489.840 ;
        RECT 504.690 489.640 505.010 489.700 ;
        RECT 570.470 489.160 570.790 489.220 ;
        RECT 876.370 489.160 876.690 489.220 ;
        RECT 570.470 489.020 876.690 489.160 ;
        RECT 570.470 488.960 570.790 489.020 ;
        RECT 876.370 488.960 876.690 489.020 ;
      LAYER via ;
        RECT 504.720 489.640 504.980 489.900 ;
        RECT 570.500 490.320 570.760 490.580 ;
        RECT 570.500 488.960 570.760 489.220 ;
        RECT 876.400 488.960 876.660 489.220 ;
      LAYER met2 ;
        RECT 504.510 500.000 504.790 504.000 ;
        RECT 504.550 498.680 504.690 500.000 ;
        RECT 504.550 498.540 504.920 498.680 ;
        RECT 504.780 489.930 504.920 498.540 ;
        RECT 570.500 490.290 570.760 490.610 ;
        RECT 504.720 489.610 504.980 489.930 ;
        RECT 570.560 489.250 570.700 490.290 ;
        RECT 570.500 488.930 570.760 489.250 ;
        RECT 876.400 488.930 876.660 489.250 ;
        RECT 876.460 82.870 876.600 488.930 ;
        RECT 876.460 82.730 877.520 82.870 ;
        RECT 877.380 2.400 877.520 82.730 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 666.150 501.400 666.470 501.460 ;
        RECT 666.150 501.260 690.070 501.400 ;
        RECT 666.150 501.200 666.470 501.260 ;
        RECT 689.930 500.380 690.070 501.260 ;
        RECT 689.930 500.240 710.770 500.380 ;
        RECT 505.840 499.700 506.160 499.760 ;
        RECT 505.840 499.560 506.990 499.700 ;
        RECT 505.840 499.500 506.160 499.560 ;
        RECT 506.850 497.720 506.990 499.560 ;
        RECT 710.630 498.340 710.770 500.240 ;
        RECT 890.170 498.340 890.490 498.400 ;
        RECT 710.630 498.200 890.490 498.340 ;
        RECT 890.170 498.140 890.490 498.200 ;
        RECT 506.530 497.520 506.990 497.720 ;
        RECT 506.530 497.460 506.850 497.520 ;
        RECT 539.650 490.860 539.970 490.920 ;
        RECT 539.650 490.720 579.670 490.860 ;
        RECT 539.650 490.660 539.970 490.720 ;
        RECT 579.530 489.840 579.670 490.720 ;
        RECT 666.150 490.180 666.470 490.240 ;
        RECT 618.400 490.040 666.470 490.180 ;
        RECT 618.400 489.840 618.540 490.040 ;
        RECT 666.150 489.980 666.470 490.040 ;
        RECT 579.530 489.700 618.540 489.840 ;
        RECT 506.530 489.500 506.850 489.560 ;
        RECT 539.650 489.500 539.970 489.560 ;
        RECT 506.530 489.360 539.970 489.500 ;
        RECT 506.530 489.300 506.850 489.360 ;
        RECT 539.650 489.300 539.970 489.360 ;
      LAYER via ;
        RECT 666.180 501.200 666.440 501.460 ;
        RECT 505.870 499.500 506.130 499.760 ;
        RECT 890.200 498.140 890.460 498.400 ;
        RECT 506.560 497.460 506.820 497.720 ;
        RECT 539.680 490.660 539.940 490.920 ;
        RECT 666.180 489.980 666.440 490.240 ;
        RECT 506.560 489.300 506.820 489.560 ;
        RECT 539.680 489.300 539.940 489.560 ;
      LAYER met2 ;
        RECT 505.890 500.000 506.170 504.000 ;
        RECT 666.180 501.170 666.440 501.490 ;
        RECT 505.930 499.790 506.070 500.000 ;
        RECT 505.870 499.470 506.130 499.790 ;
        RECT 506.560 497.430 506.820 497.750 ;
        RECT 506.620 489.590 506.760 497.430 ;
        RECT 539.680 490.630 539.940 490.950 ;
        RECT 539.740 489.590 539.880 490.630 ;
        RECT 666.240 490.270 666.380 501.170 ;
        RECT 890.200 498.110 890.460 498.430 ;
        RECT 666.180 489.950 666.440 490.270 ;
        RECT 506.560 489.270 506.820 489.590 ;
        RECT 539.680 489.270 539.940 489.590 ;
        RECT 890.260 82.870 890.400 498.110 ;
        RECT 890.260 82.730 893.160 82.870 ;
        RECT 893.020 1.770 893.160 82.730 ;
        RECT 895.110 1.770 895.670 2.400 ;
        RECT 893.020 1.630 895.670 1.770 ;
        RECT 895.110 -4.800 895.670 1.630 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 663.390 498.000 663.710 498.060 ;
        RECT 910.870 498.000 911.190 498.060 ;
        RECT 663.390 497.860 911.190 498.000 ;
        RECT 663.390 497.800 663.710 497.860 ;
        RECT 910.870 497.800 911.190 497.860 ;
        RECT 632.570 490.520 632.890 490.580 ;
        RECT 663.390 490.520 663.710 490.580 ;
        RECT 632.570 490.380 663.710 490.520 ;
        RECT 632.570 490.320 632.890 490.380 ;
        RECT 663.390 490.320 663.710 490.380 ;
        RECT 618.770 489.840 619.090 489.900 ;
        RECT 632.570 489.840 632.890 489.900 ;
        RECT 618.770 489.700 632.890 489.840 ;
        RECT 618.770 489.640 619.090 489.700 ;
        RECT 632.570 489.640 632.890 489.700 ;
        RECT 508.370 488.820 508.690 488.880 ;
        RECT 508.370 488.680 526.540 488.820 ;
        RECT 508.370 488.620 508.690 488.680 ;
        RECT 526.400 488.480 526.540 488.680 ;
        RECT 618.770 488.480 619.090 488.540 ;
        RECT 526.400 488.340 544.250 488.480 ;
        RECT 544.110 488.140 544.250 488.340 ;
        RECT 545.030 488.340 619.090 488.480 ;
        RECT 545.030 488.140 545.170 488.340 ;
        RECT 618.770 488.280 619.090 488.340 ;
        RECT 544.110 488.000 545.170 488.140 ;
      LAYER via ;
        RECT 663.420 497.800 663.680 498.060 ;
        RECT 910.900 497.800 911.160 498.060 ;
        RECT 632.600 490.320 632.860 490.580 ;
        RECT 663.420 490.320 663.680 490.580 ;
        RECT 618.800 489.640 619.060 489.900 ;
        RECT 632.600 489.640 632.860 489.900 ;
        RECT 508.400 488.620 508.660 488.880 ;
        RECT 618.800 488.280 619.060 488.540 ;
      LAYER met2 ;
        RECT 507.270 500.000 507.550 504.000 ;
        RECT 507.310 498.680 507.450 500.000 ;
        RECT 507.310 498.540 508.140 498.680 ;
        RECT 508.000 492.050 508.140 498.540 ;
        RECT 663.420 497.770 663.680 498.090 ;
        RECT 910.900 497.770 911.160 498.090 ;
        RECT 508.000 491.910 508.600 492.050 ;
        RECT 508.460 488.910 508.600 491.910 ;
        RECT 663.480 490.610 663.620 497.770 ;
        RECT 632.600 490.290 632.860 490.610 ;
        RECT 663.420 490.290 663.680 490.610 ;
        RECT 632.660 489.930 632.800 490.290 ;
        RECT 618.800 489.610 619.060 489.930 ;
        RECT 632.600 489.610 632.860 489.930 ;
        RECT 508.400 488.590 508.660 488.910 ;
        RECT 618.860 488.570 619.000 489.610 ;
        RECT 618.800 488.250 619.060 488.570 ;
        RECT 910.960 1.770 911.100 497.770 ;
        RECT 912.590 1.770 913.150 2.400 ;
        RECT 910.960 1.630 913.150 1.770 ;
        RECT 912.590 -4.800 913.150 1.630 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.690 471.140 505.010 471.200 ;
        RECT 508.830 471.140 509.150 471.200 ;
        RECT 504.690 471.000 509.150 471.140 ;
        RECT 504.690 470.940 505.010 471.000 ;
        RECT 508.830 470.940 509.150 471.000 ;
        RECT 504.690 54.300 505.010 54.360 ;
        RECT 930.650 54.300 930.970 54.360 ;
        RECT 504.690 54.160 930.970 54.300 ;
        RECT 504.690 54.100 505.010 54.160 ;
        RECT 930.650 54.100 930.970 54.160 ;
      LAYER via ;
        RECT 504.720 470.940 504.980 471.200 ;
        RECT 508.860 470.940 509.120 471.200 ;
        RECT 504.720 54.100 504.980 54.360 ;
        RECT 930.680 54.100 930.940 54.360 ;
      LAYER met2 ;
        RECT 508.650 500.000 508.930 504.000 ;
        RECT 508.690 499.020 508.830 500.000 ;
        RECT 508.690 498.880 509.060 499.020 ;
        RECT 508.920 471.230 509.060 498.880 ;
        RECT 504.720 470.910 504.980 471.230 ;
        RECT 508.860 470.910 509.120 471.230 ;
        RECT 504.780 54.390 504.920 470.910 ;
        RECT 504.720 54.070 504.980 54.390 ;
        RECT 930.680 54.070 930.940 54.390 ;
        RECT 930.740 2.400 930.880 54.070 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 509.980 498.820 510.300 499.080 ;
        RECT 510.070 497.380 510.210 498.820 ;
        RECT 510.070 497.180 510.530 497.380 ;
        RECT 510.210 497.120 510.530 497.180 ;
      LAYER via ;
        RECT 510.010 498.820 510.270 499.080 ;
        RECT 510.240 497.120 510.500 497.380 ;
      LAYER met2 ;
        RECT 510.030 500.000 510.310 504.000 ;
        RECT 510.070 499.110 510.210 500.000 ;
        RECT 510.010 498.790 510.270 499.110 ;
        RECT 510.240 497.090 510.500 497.410 ;
        RECT 510.300 483.325 510.440 497.090 ;
        RECT 510.230 482.955 510.510 483.325 ;
        RECT 946.310 53.195 946.590 53.565 ;
        RECT 946.380 1.770 946.520 53.195 ;
        RECT 948.470 1.770 949.030 2.400 ;
        RECT 946.380 1.630 949.030 1.770 ;
        RECT 948.470 -4.800 949.030 1.630 ;
      LAYER via2 ;
        RECT 510.230 483.000 510.510 483.280 ;
        RECT 946.310 53.240 946.590 53.520 ;
      LAYER met3 ;
        RECT 510.205 483.300 510.535 483.305 ;
        RECT 509.950 483.290 510.535 483.300 ;
        RECT 509.750 482.990 510.535 483.290 ;
        RECT 509.950 482.980 510.535 482.990 ;
        RECT 510.205 482.975 510.535 482.980 ;
        RECT 509.950 53.530 510.330 53.540 ;
        RECT 946.285 53.530 946.615 53.545 ;
        RECT 509.950 53.230 946.615 53.530 ;
        RECT 509.950 53.220 510.330 53.230 ;
        RECT 946.285 53.215 946.615 53.230 ;
      LAYER via3 ;
        RECT 509.980 482.980 510.300 483.300 ;
        RECT 509.980 53.220 510.300 53.540 ;
      LAYER met4 ;
        RECT 509.975 482.975 510.305 483.305 ;
        RECT 509.990 53.545 510.290 482.975 ;
        RECT 509.975 53.215 510.305 53.545 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.360 499.160 511.680 499.420 ;
        RECT 511.450 498.060 511.590 499.160 ;
        RECT 511.130 497.860 511.590 498.060 ;
        RECT 511.130 497.800 511.450 497.860 ;
        RECT 511.130 53.960 511.450 54.020 ;
        RECT 966.530 53.960 966.850 54.020 ;
        RECT 511.130 53.820 966.850 53.960 ;
        RECT 511.130 53.760 511.450 53.820 ;
        RECT 966.530 53.760 966.850 53.820 ;
      LAYER via ;
        RECT 511.390 499.160 511.650 499.420 ;
        RECT 511.160 497.800 511.420 498.060 ;
        RECT 511.160 53.760 511.420 54.020 ;
        RECT 966.560 53.760 966.820 54.020 ;
      LAYER met2 ;
        RECT 511.410 500.000 511.690 504.000 ;
        RECT 511.450 499.450 511.590 500.000 ;
        RECT 511.390 499.130 511.650 499.450 ;
        RECT 511.160 497.770 511.420 498.090 ;
        RECT 511.220 54.050 511.360 497.770 ;
        RECT 511.160 53.730 511.420 54.050 ;
        RECT 966.560 53.730 966.820 54.050 ;
        RECT 966.620 17.410 966.760 53.730 ;
        RECT 966.160 17.270 966.760 17.410 ;
        RECT 966.160 2.400 966.300 17.270 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.070 496.640 414.390 496.700 ;
        RECT 414.070 496.500 420.970 496.640 ;
        RECT 414.070 496.440 414.390 496.500 ;
        RECT 420.830 496.300 420.970 496.500 ;
        RECT 420.830 496.160 448.570 496.300 ;
        RECT 448.430 495.960 448.570 496.160 ;
        RECT 486.290 495.960 486.610 496.020 ;
        RECT 448.430 495.820 486.610 495.960 ;
        RECT 486.290 495.760 486.610 495.820 ;
      LAYER via ;
        RECT 414.100 496.440 414.360 496.700 ;
        RECT 486.320 495.760 486.580 496.020 ;
      LAYER met2 ;
        RECT 418.490 796.690 418.770 800.000 ;
        RECT 414.160 796.550 418.770 796.690 ;
        RECT 414.160 496.730 414.300 796.550 ;
        RECT 418.490 796.000 418.770 796.550 ;
        RECT 486.570 500.000 486.850 504.000 ;
        RECT 486.610 498.680 486.750 500.000 ;
        RECT 486.380 498.540 486.750 498.680 ;
        RECT 414.100 496.410 414.360 496.730 ;
        RECT 486.380 496.050 486.520 498.540 ;
        RECT 486.320 495.730 486.580 496.050 ;
        RECT 486.380 490.805 486.520 495.730 ;
        RECT 486.310 490.435 486.590 490.805 ;
        RECT 646.850 18.515 647.130 18.885 ;
        RECT 646.920 2.400 647.060 18.515 ;
        RECT 646.710 -4.800 647.270 2.400 ;
      LAYER via2 ;
        RECT 486.310 490.480 486.590 490.760 ;
        RECT 646.850 18.560 647.130 18.840 ;
      LAYER met3 ;
        RECT 486.285 490.770 486.615 490.785 ;
        RECT 488.790 490.770 489.170 490.780 ;
        RECT 486.285 490.470 489.170 490.770 ;
        RECT 486.285 490.455 486.615 490.470 ;
        RECT 488.790 490.460 489.170 490.470 ;
        RECT 488.790 18.850 489.170 18.860 ;
        RECT 646.825 18.850 647.155 18.865 ;
        RECT 488.790 18.550 647.155 18.850 ;
        RECT 488.790 18.540 489.170 18.550 ;
        RECT 646.825 18.535 647.155 18.550 ;
      LAYER via3 ;
        RECT 488.820 490.460 489.140 490.780 ;
        RECT 488.820 18.540 489.140 18.860 ;
      LAYER met4 ;
        RECT 488.815 490.455 489.145 490.785 ;
        RECT 488.830 18.865 489.130 490.455 ;
        RECT 488.815 18.535 489.145 18.865 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.590 53.620 511.910 53.680 ;
        RECT 984.010 53.620 984.330 53.680 ;
        RECT 511.590 53.480 984.330 53.620 ;
        RECT 511.590 53.420 511.910 53.480 ;
        RECT 984.010 53.420 984.330 53.480 ;
      LAYER via ;
        RECT 511.620 53.420 511.880 53.680 ;
        RECT 984.040 53.420 984.300 53.680 ;
      LAYER met2 ;
        RECT 512.790 500.000 513.070 504.000 ;
        RECT 512.830 498.965 512.970 500.000 ;
        RECT 512.760 498.595 513.040 498.965 ;
        RECT 512.070 497.915 512.350 498.285 ;
        RECT 512.140 472.500 512.280 497.915 ;
        RECT 511.680 472.360 512.280 472.500 ;
        RECT 511.680 53.710 511.820 472.360 ;
        RECT 511.620 53.390 511.880 53.710 ;
        RECT 984.040 53.390 984.300 53.710 ;
        RECT 984.100 2.400 984.240 53.390 ;
        RECT 983.890 -4.800 984.450 2.400 ;
      LAYER via2 ;
        RECT 512.760 498.640 513.040 498.920 ;
        RECT 512.070 497.960 512.350 498.240 ;
      LAYER met3 ;
        RECT 512.735 498.615 513.065 498.945 ;
        RECT 512.045 498.250 512.375 498.265 ;
        RECT 512.750 498.250 513.050 498.615 ;
        RECT 512.045 497.950 513.050 498.250 ;
        RECT 512.045 497.935 512.375 497.950 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 514.120 499.160 514.440 499.420 ;
        RECT 513.430 497.660 513.750 497.720 ;
        RECT 514.210 497.660 514.350 499.160 ;
        RECT 513.430 497.520 514.350 497.660 ;
        RECT 513.430 497.460 513.750 497.520 ;
        RECT 512.050 465.360 512.370 465.420 ;
        RECT 513.430 465.360 513.750 465.420 ;
        RECT 512.050 465.220 513.750 465.360 ;
        RECT 512.050 465.160 512.370 465.220 ;
        RECT 513.430 465.160 513.750 465.220 ;
        RECT 512.050 61.100 512.370 61.160 ;
        RECT 1001.490 61.100 1001.810 61.160 ;
        RECT 512.050 60.960 1001.810 61.100 ;
        RECT 512.050 60.900 512.370 60.960 ;
        RECT 1001.490 60.900 1001.810 60.960 ;
      LAYER via ;
        RECT 514.150 499.160 514.410 499.420 ;
        RECT 513.460 497.460 513.720 497.720 ;
        RECT 512.080 465.160 512.340 465.420 ;
        RECT 513.460 465.160 513.720 465.420 ;
        RECT 512.080 60.900 512.340 61.160 ;
        RECT 1001.520 60.900 1001.780 61.160 ;
      LAYER met2 ;
        RECT 514.170 500.000 514.450 504.000 ;
        RECT 514.210 499.450 514.350 500.000 ;
        RECT 514.150 499.130 514.410 499.450 ;
        RECT 513.460 497.430 513.720 497.750 ;
        RECT 513.520 465.450 513.660 497.430 ;
        RECT 512.080 465.130 512.340 465.450 ;
        RECT 513.460 465.130 513.720 465.450 ;
        RECT 512.140 61.190 512.280 465.130 ;
        RECT 512.080 60.870 512.340 61.190 ;
        RECT 1001.520 60.870 1001.780 61.190 ;
        RECT 1001.580 2.400 1001.720 60.870 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.550 500.000 515.830 504.000 ;
        RECT 515.590 498.965 515.730 500.000 ;
        RECT 515.520 498.595 515.800 498.965 ;
        RECT 1017.150 60.675 1017.430 61.045 ;
        RECT 1017.220 1.770 1017.360 60.675 ;
        RECT 1019.310 1.770 1019.870 2.400 ;
        RECT 1017.220 1.630 1019.870 1.770 ;
        RECT 1019.310 -4.800 1019.870 1.630 ;
      LAYER via2 ;
        RECT 515.520 498.640 515.800 498.920 ;
        RECT 1017.150 60.720 1017.430 61.000 ;
      LAYER met3 ;
        RECT 515.495 498.940 515.825 498.945 ;
        RECT 515.470 498.930 515.850 498.940 ;
        RECT 515.040 498.630 515.850 498.930 ;
        RECT 515.470 498.620 515.850 498.630 ;
        RECT 515.495 498.615 515.825 498.620 ;
        RECT 515.470 61.010 515.850 61.020 ;
        RECT 1017.125 61.010 1017.455 61.025 ;
        RECT 515.470 60.710 1017.455 61.010 ;
        RECT 515.470 60.700 515.850 60.710 ;
        RECT 1017.125 60.695 1017.455 60.710 ;
      LAYER via3 ;
        RECT 515.500 498.620 515.820 498.940 ;
        RECT 515.500 60.700 515.820 61.020 ;
      LAYER met4 ;
        RECT 515.495 498.615 515.825 498.945 ;
        RECT 515.510 61.025 515.810 498.615 ;
        RECT 515.495 60.695 515.825 61.025 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.930 500.000 517.210 504.000 ;
        RECT 516.970 499.645 517.110 500.000 ;
        RECT 516.900 499.275 517.180 499.645 ;
        RECT 1035.090 59.995 1035.370 60.365 ;
        RECT 1035.160 1.770 1035.300 59.995 ;
        RECT 1036.790 1.770 1037.350 2.400 ;
        RECT 1035.160 1.630 1037.350 1.770 ;
        RECT 1036.790 -4.800 1037.350 1.630 ;
      LAYER via2 ;
        RECT 516.900 499.320 517.180 499.600 ;
        RECT 1035.090 60.040 1035.370 60.320 ;
      LAYER met3 ;
        RECT 515.470 499.610 515.850 499.620 ;
        RECT 516.875 499.610 517.205 499.625 ;
        RECT 515.470 499.310 517.205 499.610 ;
        RECT 515.470 499.300 515.850 499.310 ;
        RECT 516.875 499.295 517.205 499.310 ;
        RECT 516.390 60.330 516.770 60.340 ;
        RECT 1035.065 60.330 1035.395 60.345 ;
        RECT 516.390 60.030 1035.395 60.330 ;
        RECT 516.390 60.020 516.770 60.030 ;
        RECT 1035.065 60.015 1035.395 60.030 ;
      LAYER via3 ;
        RECT 515.500 499.300 515.820 499.620 ;
        RECT 516.420 60.020 516.740 60.340 ;
      LAYER met4 ;
        RECT 515.495 499.610 515.825 499.625 ;
        RECT 515.495 499.310 516.730 499.610 ;
        RECT 515.495 499.295 515.825 499.310 ;
        RECT 516.430 60.345 516.730 499.310 ;
        RECT 516.415 60.015 516.745 60.345 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.570 19.280 517.890 19.340 ;
        RECT 1054.850 19.280 1055.170 19.340 ;
        RECT 517.570 19.140 1055.170 19.280 ;
        RECT 517.570 19.080 517.890 19.140 ;
        RECT 1054.850 19.080 1055.170 19.140 ;
      LAYER via ;
        RECT 517.600 19.080 517.860 19.340 ;
        RECT 1054.880 19.080 1055.140 19.340 ;
      LAYER met2 ;
        RECT 518.310 500.000 518.590 504.000 ;
        RECT 518.350 499.020 518.490 500.000 ;
        RECT 518.120 498.880 518.490 499.020 ;
        RECT 518.120 492.560 518.260 498.880 ;
        RECT 517.660 492.420 518.260 492.560 ;
        RECT 517.660 19.370 517.800 492.420 ;
        RECT 517.600 19.050 517.860 19.370 ;
        RECT 1054.880 19.050 1055.140 19.370 ;
        RECT 1054.940 2.400 1055.080 19.050 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 519.640 499.500 519.960 499.760 ;
        RECT 519.730 498.000 519.870 499.500 ;
        RECT 519.730 497.860 521.020 498.000 ;
        RECT 519.410 496.980 519.730 497.040 ;
        RECT 520.880 496.980 521.020 497.860 ;
        RECT 519.410 496.840 521.020 496.980 ;
        RECT 519.410 496.780 519.730 496.840 ;
        RECT 519.410 60.760 519.730 60.820 ;
        RECT 1072.330 60.760 1072.650 60.820 ;
        RECT 519.410 60.620 1072.650 60.760 ;
        RECT 519.410 60.560 519.730 60.620 ;
        RECT 1072.330 60.560 1072.650 60.620 ;
      LAYER via ;
        RECT 519.670 499.500 519.930 499.760 ;
        RECT 519.440 496.780 519.700 497.040 ;
        RECT 519.440 60.560 519.700 60.820 ;
        RECT 1072.360 60.560 1072.620 60.820 ;
      LAYER met2 ;
        RECT 519.690 500.000 519.970 504.000 ;
        RECT 519.730 499.790 519.870 500.000 ;
        RECT 519.670 499.470 519.930 499.790 ;
        RECT 519.440 496.750 519.700 497.070 ;
        RECT 519.500 60.850 519.640 496.750 ;
        RECT 519.440 60.530 519.700 60.850 ;
        RECT 1072.360 60.530 1072.620 60.850 ;
        RECT 1072.420 2.400 1072.560 60.530 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 519.870 60.420 520.190 60.480 ;
        RECT 1090.730 60.420 1091.050 60.480 ;
        RECT 519.870 60.280 1091.050 60.420 ;
        RECT 519.870 60.220 520.190 60.280 ;
        RECT 1090.730 60.220 1091.050 60.280 ;
      LAYER via ;
        RECT 519.900 60.220 520.160 60.480 ;
        RECT 1090.760 60.220 1091.020 60.480 ;
      LAYER met2 ;
        RECT 521.070 500.000 521.350 504.000 ;
        RECT 521.110 499.645 521.250 500.000 ;
        RECT 521.040 499.275 521.320 499.645 ;
        RECT 519.890 497.235 520.170 497.605 ;
        RECT 519.960 60.510 520.100 497.235 ;
        RECT 519.900 60.190 520.160 60.510 ;
        RECT 1090.760 60.190 1091.020 60.510 ;
        RECT 1090.820 34.570 1090.960 60.190 ;
        RECT 1090.360 34.430 1090.960 34.570 ;
        RECT 1090.360 2.400 1090.500 34.430 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
      LAYER via2 ;
        RECT 521.040 499.320 521.320 499.600 ;
        RECT 519.890 497.280 520.170 497.560 ;
      LAYER met3 ;
        RECT 521.015 499.610 521.345 499.625 ;
        RECT 519.880 499.310 521.345 499.610 ;
        RECT 519.880 497.585 520.180 499.310 ;
        RECT 521.015 499.295 521.345 499.310 ;
        RECT 519.865 497.255 520.195 497.585 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.450 500.000 522.730 504.000 ;
        RECT 522.490 499.815 522.630 500.000 ;
        RECT 522.420 499.445 522.700 499.815 ;
        RECT 1105.470 66.795 1105.750 67.165 ;
        RECT 1105.540 1.770 1105.680 66.795 ;
        RECT 1107.630 1.770 1108.190 2.400 ;
        RECT 1105.540 1.630 1108.190 1.770 ;
        RECT 1107.630 -4.800 1108.190 1.630 ;
      LAYER via2 ;
        RECT 522.420 499.490 522.700 499.770 ;
        RECT 1105.470 66.840 1105.750 67.120 ;
      LAYER met3 ;
        RECT 522.395 499.780 522.725 499.795 ;
        RECT 522.180 499.620 522.725 499.780 ;
        RECT 521.910 499.465 522.725 499.620 ;
        RECT 521.910 499.310 522.480 499.465 ;
        RECT 521.910 499.300 522.290 499.310 ;
        RECT 521.910 67.130 522.290 67.140 ;
        RECT 1105.445 67.130 1105.775 67.145 ;
        RECT 521.910 66.830 1105.775 67.130 ;
        RECT 521.910 66.820 522.290 66.830 ;
        RECT 1105.445 66.815 1105.775 66.830 ;
      LAYER via3 ;
        RECT 521.940 499.300 522.260 499.620 ;
        RECT 521.940 66.820 522.260 67.140 ;
      LAYER met4 ;
        RECT 521.935 499.295 522.265 499.625 ;
        RECT 521.950 67.145 522.250 499.295 ;
        RECT 521.935 66.815 522.265 67.145 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.830 500.000 524.110 504.000 ;
        RECT 523.870 499.815 524.010 500.000 ;
        RECT 523.800 499.445 524.080 499.815 ;
        RECT 1125.710 66.115 1125.990 66.485 ;
        RECT 1125.780 2.400 1125.920 66.115 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
      LAYER via2 ;
        RECT 523.800 499.490 524.080 499.770 ;
        RECT 1125.710 66.160 1125.990 66.440 ;
      LAYER met3 ;
        RECT 523.775 499.620 524.105 499.795 ;
        RECT 523.750 499.610 524.130 499.620 ;
        RECT 523.750 499.310 524.390 499.610 ;
        RECT 523.750 499.300 524.130 499.310 ;
        RECT 522.830 66.450 523.210 66.460 ;
        RECT 1125.685 66.450 1126.015 66.465 ;
        RECT 522.830 66.150 1126.015 66.450 ;
        RECT 522.830 66.140 523.210 66.150 ;
        RECT 1125.685 66.135 1126.015 66.150 ;
      LAYER via3 ;
        RECT 523.780 499.300 524.100 499.620 ;
        RECT 522.860 66.140 523.180 66.460 ;
      LAYER met4 ;
        RECT 523.775 499.610 524.105 499.625 ;
        RECT 522.870 499.310 524.105 499.610 ;
        RECT 522.870 66.465 523.170 499.310 ;
        RECT 523.775 499.295 524.105 499.310 ;
        RECT 522.855 66.135 523.185 66.465 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.930 492.220 525.250 492.280 ;
        RECT 1138.570 492.220 1138.890 492.280 ;
        RECT 524.930 492.080 1138.890 492.220 ;
        RECT 524.930 492.020 525.250 492.080 ;
        RECT 1138.570 492.020 1138.890 492.080 ;
      LAYER via ;
        RECT 524.960 492.020 525.220 492.280 ;
        RECT 1138.600 492.020 1138.860 492.280 ;
      LAYER met2 ;
        RECT 525.210 500.000 525.490 504.000 ;
        RECT 525.250 498.850 525.390 500.000 ;
        RECT 525.020 498.710 525.390 498.850 ;
        RECT 525.020 492.310 525.160 498.710 ;
        RECT 524.960 491.990 525.220 492.310 ;
        RECT 1138.600 491.990 1138.860 492.310 ;
        RECT 1138.660 82.870 1138.800 491.990 ;
        RECT 1138.660 82.730 1141.560 82.870 ;
        RECT 1141.420 1.770 1141.560 82.730 ;
        RECT 1143.510 1.770 1144.070 2.400 ;
        RECT 1141.420 1.630 1144.070 1.770 ;
        RECT 1143.510 -4.800 1144.070 1.630 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 487.900 499.500 488.220 499.760 ;
        RECT 487.990 498.400 488.130 499.500 ;
        RECT 487.990 498.200 488.450 498.400 ;
        RECT 488.130 498.140 488.450 498.200 ;
        RECT 488.590 18.600 488.910 18.660 ;
        RECT 664.770 18.600 665.090 18.660 ;
        RECT 488.590 18.460 665.090 18.600 ;
        RECT 488.590 18.400 488.910 18.460 ;
        RECT 664.770 18.400 665.090 18.460 ;
      LAYER via ;
        RECT 487.930 499.500 488.190 499.760 ;
        RECT 488.160 498.140 488.420 498.400 ;
        RECT 488.620 18.400 488.880 18.660 ;
        RECT 664.800 18.400 665.060 18.660 ;
      LAYER met2 ;
        RECT 487.950 500.000 488.230 504.000 ;
        RECT 487.990 499.790 488.130 500.000 ;
        RECT 487.930 499.470 488.190 499.790 ;
        RECT 488.160 498.110 488.420 498.430 ;
        RECT 488.220 476.170 488.360 498.110 ;
        RECT 487.760 476.030 488.360 476.170 ;
        RECT 487.760 448.570 487.900 476.030 ;
        RECT 487.760 448.430 488.820 448.570 ;
        RECT 488.680 18.690 488.820 448.430 ;
        RECT 488.620 18.370 488.880 18.690 ;
        RECT 664.800 18.370 665.060 18.690 ;
        RECT 664.860 2.400 665.000 18.370 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 526.540 498.820 526.860 499.080 ;
        RECT 526.630 497.720 526.770 498.820 ;
        RECT 526.630 497.520 527.090 497.720 ;
        RECT 526.770 497.460 527.090 497.520 ;
        RECT 526.770 492.560 527.090 492.620 ;
        RECT 1159.270 492.560 1159.590 492.620 ;
        RECT 526.770 492.420 1159.590 492.560 ;
        RECT 526.770 492.360 527.090 492.420 ;
        RECT 1159.270 492.360 1159.590 492.420 ;
      LAYER via ;
        RECT 526.570 498.820 526.830 499.080 ;
        RECT 526.800 497.460 527.060 497.720 ;
        RECT 526.800 492.360 527.060 492.620 ;
        RECT 1159.300 492.360 1159.560 492.620 ;
      LAYER met2 ;
        RECT 526.590 500.000 526.870 504.000 ;
        RECT 526.630 499.110 526.770 500.000 ;
        RECT 526.570 498.790 526.830 499.110 ;
        RECT 526.800 497.430 527.060 497.750 ;
        RECT 526.860 492.650 527.000 497.430 ;
        RECT 526.800 492.330 527.060 492.650 ;
        RECT 1159.300 492.330 1159.560 492.650 ;
        RECT 1159.360 1.770 1159.500 492.330 ;
        RECT 1160.990 1.770 1161.550 2.400 ;
        RECT 1159.360 1.630 1161.550 1.770 ;
        RECT 1160.990 -4.800 1161.550 1.630 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 526.310 74.700 526.630 74.760 ;
        RECT 1179.050 74.700 1179.370 74.760 ;
        RECT 526.310 74.560 1179.370 74.700 ;
        RECT 526.310 74.500 526.630 74.560 ;
        RECT 1179.050 74.500 1179.370 74.560 ;
      LAYER via ;
        RECT 526.340 74.500 526.600 74.760 ;
        RECT 1179.080 74.500 1179.340 74.760 ;
      LAYER met2 ;
        RECT 527.970 500.000 528.250 504.000 ;
        RECT 528.010 498.965 528.150 500.000 ;
        RECT 527.940 498.595 528.220 498.965 ;
        RECT 526.330 491.795 526.610 492.165 ;
        RECT 526.400 74.790 526.540 491.795 ;
        RECT 526.340 74.470 526.600 74.790 ;
        RECT 1179.080 74.470 1179.340 74.790 ;
        RECT 1179.140 2.400 1179.280 74.470 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
      LAYER via2 ;
        RECT 527.940 498.640 528.220 498.920 ;
        RECT 526.330 491.840 526.610 492.120 ;
      LAYER met3 ;
        RECT 526.510 498.930 526.890 498.940 ;
        RECT 527.915 498.930 528.245 498.945 ;
        RECT 526.510 498.630 528.245 498.930 ;
        RECT 526.510 498.620 526.890 498.630 ;
        RECT 527.915 498.615 528.245 498.630 ;
        RECT 526.305 492.140 526.635 492.145 ;
        RECT 526.305 492.130 526.890 492.140 ;
        RECT 526.080 491.830 526.890 492.130 ;
        RECT 526.305 491.820 526.890 491.830 ;
        RECT 526.305 491.815 526.635 491.820 ;
      LAYER via3 ;
        RECT 526.540 498.620 526.860 498.940 ;
        RECT 526.540 491.820 526.860 492.140 ;
      LAYER met4 ;
        RECT 526.535 498.615 526.865 498.945 ;
        RECT 526.550 492.145 526.850 498.615 ;
        RECT 526.535 491.815 526.865 492.145 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 529.300 499.360 529.620 499.420 ;
        RECT 529.300 499.160 529.760 499.360 ;
        RECT 529.620 498.400 529.760 499.160 ;
        RECT 529.530 498.140 529.850 498.400 ;
        RECT 524.470 483.040 524.790 483.100 ;
        RECT 529.530 483.040 529.850 483.100 ;
        RECT 524.470 482.900 529.850 483.040 ;
        RECT 524.470 482.840 524.790 482.900 ;
        RECT 529.530 482.840 529.850 482.900 ;
        RECT 524.470 33.900 524.790 33.960 ;
        RECT 1196.530 33.900 1196.850 33.960 ;
        RECT 524.470 33.760 1196.850 33.900 ;
        RECT 524.470 33.700 524.790 33.760 ;
        RECT 1196.530 33.700 1196.850 33.760 ;
      LAYER via ;
        RECT 529.330 499.160 529.590 499.420 ;
        RECT 529.560 498.140 529.820 498.400 ;
        RECT 524.500 482.840 524.760 483.100 ;
        RECT 529.560 482.840 529.820 483.100 ;
        RECT 524.500 33.700 524.760 33.960 ;
        RECT 1196.560 33.700 1196.820 33.960 ;
      LAYER met2 ;
        RECT 529.350 500.000 529.630 504.000 ;
        RECT 529.390 499.450 529.530 500.000 ;
        RECT 529.330 499.130 529.590 499.450 ;
        RECT 529.560 498.110 529.820 498.430 ;
        RECT 529.620 483.130 529.760 498.110 ;
        RECT 524.500 482.810 524.760 483.130 ;
        RECT 529.560 482.810 529.820 483.130 ;
        RECT 524.560 33.990 524.700 482.810 ;
        RECT 524.500 33.670 524.760 33.990 ;
        RECT 1196.560 33.670 1196.820 33.990 ;
        RECT 1196.620 2.400 1196.760 33.670 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 530.680 499.500 531.000 499.760 ;
        RECT 530.770 499.080 530.910 499.500 ;
        RECT 530.450 498.880 530.910 499.080 ;
        RECT 530.450 498.820 530.770 498.880 ;
      LAYER via ;
        RECT 530.710 499.500 530.970 499.760 ;
        RECT 530.480 498.820 530.740 499.080 ;
      LAYER met2 ;
        RECT 530.730 500.000 531.010 504.000 ;
        RECT 530.770 499.790 530.910 500.000 ;
        RECT 530.710 499.470 530.970 499.790 ;
        RECT 530.480 498.790 530.740 499.110 ;
        RECT 530.540 488.085 530.680 498.790 ;
        RECT 530.470 487.715 530.750 488.085 ;
        RECT 1214.950 75.635 1215.230 76.005 ;
        RECT 1215.020 34.570 1215.160 75.635 ;
        RECT 1214.560 34.430 1215.160 34.570 ;
        RECT 1214.560 2.400 1214.700 34.430 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
      LAYER via2 ;
        RECT 530.470 487.760 530.750 488.040 ;
        RECT 1214.950 75.680 1215.230 75.960 ;
      LAYER met3 ;
        RECT 530.445 488.060 530.775 488.065 ;
        RECT 530.190 488.050 530.775 488.060 ;
        RECT 529.990 487.750 530.775 488.050 ;
        RECT 530.190 487.740 530.775 487.750 ;
        RECT 530.445 487.735 530.775 487.740 ;
        RECT 530.190 75.970 530.570 75.980 ;
        RECT 1214.925 75.970 1215.255 75.985 ;
        RECT 530.190 75.670 1215.255 75.970 ;
        RECT 530.190 75.660 530.570 75.670 ;
        RECT 1214.925 75.655 1215.255 75.670 ;
      LAYER via3 ;
        RECT 530.220 487.740 530.540 488.060 ;
        RECT 530.220 75.660 530.540 75.980 ;
      LAYER met4 ;
        RECT 530.215 487.735 530.545 488.065 ;
        RECT 530.230 75.985 530.530 487.735 ;
        RECT 530.215 75.655 530.545 75.985 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 532.060 499.500 532.380 499.760 ;
        RECT 532.150 497.320 532.290 499.500 ;
        RECT 536.430 497.320 536.750 497.380 ;
        RECT 532.150 497.180 536.750 497.320 ;
        RECT 536.430 497.120 536.750 497.180 ;
        RECT 536.430 18.940 536.750 19.000 ;
        RECT 1231.950 18.940 1232.270 19.000 ;
        RECT 536.430 18.800 1232.270 18.940 ;
        RECT 536.430 18.740 536.750 18.800 ;
        RECT 1231.950 18.740 1232.270 18.800 ;
      LAYER via ;
        RECT 532.090 499.500 532.350 499.760 ;
        RECT 536.460 497.120 536.720 497.380 ;
        RECT 536.460 18.740 536.720 19.000 ;
        RECT 1231.980 18.740 1232.240 19.000 ;
      LAYER met2 ;
        RECT 532.110 500.000 532.390 504.000 ;
        RECT 532.150 499.790 532.290 500.000 ;
        RECT 532.090 499.470 532.350 499.790 ;
        RECT 536.460 497.090 536.720 497.410 ;
        RECT 536.520 19.030 536.660 497.090 ;
        RECT 536.460 18.710 536.720 19.030 ;
        RECT 1231.980 18.710 1232.240 19.030 ;
        RECT 1232.040 2.400 1232.180 18.710 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 533.670 74.360 533.990 74.420 ;
        RECT 1249.890 74.360 1250.210 74.420 ;
        RECT 533.670 74.220 1250.210 74.360 ;
        RECT 533.670 74.160 533.990 74.220 ;
        RECT 1249.890 74.160 1250.210 74.220 ;
      LAYER via ;
        RECT 533.700 74.160 533.960 74.420 ;
        RECT 1249.920 74.160 1250.180 74.420 ;
      LAYER met2 ;
        RECT 533.490 500.000 533.770 504.000 ;
        RECT 533.530 498.680 533.670 500.000 ;
        RECT 533.530 498.540 533.900 498.680 ;
        RECT 533.760 74.450 533.900 498.540 ;
        RECT 533.700 74.130 533.960 74.450 ;
        RECT 1249.920 74.130 1250.180 74.450 ;
        RECT 1249.980 2.400 1250.120 74.130 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 534.820 499.500 535.140 499.760 ;
        RECT 534.130 497.660 534.450 497.720 ;
        RECT 534.910 497.660 535.050 499.500 ;
        RECT 534.130 497.520 535.050 497.660 ;
        RECT 534.130 497.460 534.450 497.520 ;
        RECT 533.210 482.700 533.530 482.760 ;
        RECT 534.130 482.700 534.450 482.760 ;
        RECT 533.210 482.560 534.450 482.700 ;
        RECT 533.210 482.500 533.530 482.560 ;
        RECT 534.130 482.500 534.450 482.560 ;
        RECT 533.210 74.020 533.530 74.080 ;
        RECT 1267.370 74.020 1267.690 74.080 ;
        RECT 533.210 73.880 1267.690 74.020 ;
        RECT 533.210 73.820 533.530 73.880 ;
        RECT 1267.370 73.820 1267.690 73.880 ;
      LAYER via ;
        RECT 534.850 499.500 535.110 499.760 ;
        RECT 534.160 497.460 534.420 497.720 ;
        RECT 533.240 482.500 533.500 482.760 ;
        RECT 534.160 482.500 534.420 482.760 ;
        RECT 533.240 73.820 533.500 74.080 ;
        RECT 1267.400 73.820 1267.660 74.080 ;
      LAYER met2 ;
        RECT 534.870 500.000 535.150 504.000 ;
        RECT 534.910 499.790 535.050 500.000 ;
        RECT 534.850 499.470 535.110 499.790 ;
        RECT 534.160 497.430 534.420 497.750 ;
        RECT 534.220 482.790 534.360 497.430 ;
        RECT 533.240 482.470 533.500 482.790 ;
        RECT 534.160 482.470 534.420 482.790 ;
        RECT 533.300 74.110 533.440 482.470 ;
        RECT 533.240 73.790 533.500 74.110 ;
        RECT 1267.400 73.790 1267.660 74.110 ;
        RECT 1267.460 2.400 1267.600 73.790 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 536.200 499.500 536.520 499.760 ;
        RECT 536.290 498.680 536.430 499.500 ;
        RECT 536.290 498.540 537.120 498.680 ;
        RECT 536.980 498.400 537.120 498.540 ;
        RECT 536.890 498.140 537.210 498.400 ;
      LAYER via ;
        RECT 536.230 499.500 536.490 499.760 ;
        RECT 536.920 498.140 537.180 498.400 ;
      LAYER met2 ;
        RECT 536.250 500.000 536.530 504.000 ;
        RECT 536.290 499.790 536.430 500.000 ;
        RECT 536.230 499.470 536.490 499.790 ;
        RECT 536.920 498.110 537.180 498.430 ;
        RECT 536.980 491.485 537.120 498.110 ;
        RECT 536.910 491.115 537.190 491.485 ;
        RECT 1283.490 74.955 1283.770 75.325 ;
        RECT 1283.560 1.770 1283.700 74.955 ;
        RECT 1285.190 1.770 1285.750 2.400 ;
        RECT 1283.560 1.630 1285.750 1.770 ;
        RECT 1285.190 -4.800 1285.750 1.630 ;
      LAYER via2 ;
        RECT 536.910 491.160 537.190 491.440 ;
        RECT 1283.490 75.000 1283.770 75.280 ;
      LAYER met3 ;
        RECT 535.710 491.450 536.090 491.460 ;
        RECT 536.885 491.450 537.215 491.465 ;
        RECT 535.710 491.150 537.215 491.450 ;
        RECT 535.710 491.140 536.090 491.150 ;
        RECT 536.885 491.135 537.215 491.150 ;
        RECT 535.710 75.290 536.090 75.300 ;
        RECT 1283.465 75.290 1283.795 75.305 ;
        RECT 535.710 74.990 1283.795 75.290 ;
        RECT 535.710 74.980 536.090 74.990 ;
        RECT 1283.465 74.975 1283.795 74.990 ;
      LAYER via3 ;
        RECT 535.740 491.140 536.060 491.460 ;
        RECT 535.740 74.980 536.060 75.300 ;
      LAYER met4 ;
        RECT 535.735 491.135 536.065 491.465 ;
        RECT 535.750 75.305 536.050 491.135 ;
        RECT 535.735 74.975 536.065 75.305 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.630 500.000 537.910 504.000 ;
        RECT 537.670 499.020 537.810 500.000 ;
        RECT 537.670 498.965 538.040 499.020 ;
        RECT 537.670 498.880 538.110 498.965 ;
        RECT 537.830 498.595 538.110 498.880 ;
        RECT 1303.270 38.235 1303.550 38.605 ;
        RECT 1303.340 2.400 1303.480 38.235 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
      LAYER via2 ;
        RECT 537.830 498.640 538.110 498.920 ;
        RECT 1303.270 38.280 1303.550 38.560 ;
      LAYER met3 ;
        RECT 537.805 498.615 538.135 498.945 ;
        RECT 537.820 498.260 538.120 498.615 ;
        RECT 537.550 497.950 538.120 498.260 ;
        RECT 537.550 497.940 537.930 497.950 ;
        RECT 537.550 38.570 537.930 38.580 ;
        RECT 1303.245 38.570 1303.575 38.585 ;
        RECT 537.550 38.270 1303.575 38.570 ;
        RECT 537.550 38.260 537.930 38.270 ;
        RECT 1303.245 38.255 1303.575 38.270 ;
      LAYER via3 ;
        RECT 537.580 497.940 537.900 498.260 ;
        RECT 537.580 38.260 537.900 38.580 ;
      LAYER met4 ;
        RECT 537.575 497.935 537.905 498.265 ;
        RECT 537.590 38.585 537.890 497.935 ;
        RECT 537.575 38.255 537.905 38.585 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 539.050 499.900 543.790 500.040 ;
        RECT 539.050 499.760 539.190 499.900 ;
        RECT 538.960 499.500 539.280 499.760 ;
        RECT 543.650 498.740 543.790 499.900 ;
        RECT 543.650 498.540 544.110 498.740 ;
        RECT 543.790 498.480 544.110 498.540 ;
        RECT 543.790 492.900 544.110 492.960 ;
        RECT 1317.970 492.900 1318.290 492.960 ;
        RECT 543.790 492.760 1318.290 492.900 ;
        RECT 543.790 492.700 544.110 492.760 ;
        RECT 1317.970 492.700 1318.290 492.760 ;
      LAYER via ;
        RECT 538.990 499.500 539.250 499.760 ;
        RECT 543.820 498.480 544.080 498.740 ;
        RECT 543.820 492.700 544.080 492.960 ;
        RECT 1318.000 492.700 1318.260 492.960 ;
      LAYER met2 ;
        RECT 539.010 500.000 539.290 504.000 ;
        RECT 539.050 499.790 539.190 500.000 ;
        RECT 538.990 499.470 539.250 499.790 ;
        RECT 543.820 498.450 544.080 498.770 ;
        RECT 543.880 492.990 544.020 498.450 ;
        RECT 543.820 492.670 544.080 492.990 ;
        RECT 1318.000 492.670 1318.260 492.990 ;
        RECT 1318.060 82.870 1318.200 492.670 ;
        RECT 1318.060 82.730 1320.960 82.870 ;
        RECT 1320.820 2.400 1320.960 82.730 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 489.050 486.440 489.370 486.500 ;
        RECT 489.050 486.300 616.700 486.440 ;
        RECT 489.050 486.240 489.370 486.300 ;
        RECT 616.560 486.100 616.700 486.300 ;
        RECT 639.010 486.100 639.330 486.160 ;
        RECT 616.560 485.960 639.330 486.100 ;
        RECT 639.010 485.900 639.330 485.960 ;
        RECT 640.390 19.960 640.710 20.020 ;
        RECT 682.250 19.960 682.570 20.020 ;
        RECT 640.390 19.820 682.570 19.960 ;
        RECT 640.390 19.760 640.710 19.820 ;
        RECT 682.250 19.760 682.570 19.820 ;
      LAYER via ;
        RECT 489.080 486.240 489.340 486.500 ;
        RECT 639.040 485.900 639.300 486.160 ;
        RECT 640.420 19.760 640.680 20.020 ;
        RECT 682.280 19.760 682.540 20.020 ;
      LAYER met2 ;
        RECT 489.330 500.000 489.610 504.000 ;
        RECT 489.370 498.850 489.510 500.000 ;
        RECT 489.140 498.710 489.510 498.850 ;
        RECT 489.140 486.530 489.280 498.710 ;
        RECT 489.080 486.210 489.340 486.530 ;
        RECT 639.040 485.870 639.300 486.190 ;
        RECT 639.100 448.570 639.240 485.870 ;
        RECT 639.100 448.430 640.620 448.570 ;
        RECT 640.480 20.050 640.620 448.430 ;
        RECT 640.420 19.730 640.680 20.050 ;
        RECT 682.280 19.730 682.540 20.050 ;
        RECT 682.340 2.400 682.480 19.730 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 540.340 499.700 540.660 499.760 ;
        RECT 539.970 499.560 540.660 499.700 ;
        RECT 539.970 499.020 540.110 499.560 ;
        RECT 540.340 499.500 540.660 499.560 ;
        RECT 539.970 498.880 540.340 499.020 ;
        RECT 540.200 498.400 540.340 498.880 ;
        RECT 540.110 498.140 540.430 498.400 ;
        RECT 540.110 81.160 540.430 81.220 ;
        RECT 1338.670 81.160 1338.990 81.220 ;
        RECT 540.110 81.020 1338.990 81.160 ;
        RECT 540.110 80.960 540.430 81.020 ;
        RECT 1338.670 80.960 1338.990 81.020 ;
      LAYER via ;
        RECT 540.370 499.500 540.630 499.760 ;
        RECT 540.140 498.140 540.400 498.400 ;
        RECT 540.140 80.960 540.400 81.220 ;
        RECT 1338.700 80.960 1338.960 81.220 ;
      LAYER met2 ;
        RECT 540.390 500.000 540.670 504.000 ;
        RECT 540.430 499.790 540.570 500.000 ;
        RECT 540.370 499.470 540.630 499.790 ;
        RECT 540.140 498.110 540.400 498.430 ;
        RECT 540.200 81.250 540.340 498.110 ;
        RECT 540.140 80.930 540.400 81.250 ;
        RECT 1338.700 80.930 1338.960 81.250 ;
        RECT 1338.760 2.400 1338.900 80.930 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 541.720 499.160 542.040 499.420 ;
        RECT 541.810 498.000 541.950 499.160 ;
        RECT 542.870 498.000 543.190 498.060 ;
        RECT 541.810 497.860 543.190 498.000 ;
        RECT 542.870 497.800 543.190 497.860 ;
        RECT 540.570 471.820 540.890 471.880 ;
        RECT 542.410 471.820 542.730 471.880 ;
        RECT 540.570 471.680 542.730 471.820 ;
        RECT 540.570 471.620 540.890 471.680 ;
        RECT 542.410 471.620 542.730 471.680 ;
        RECT 540.570 80.820 540.890 80.880 ;
        RECT 1353.850 80.820 1354.170 80.880 ;
        RECT 540.570 80.680 1354.170 80.820 ;
        RECT 540.570 80.620 540.890 80.680 ;
        RECT 1353.850 80.620 1354.170 80.680 ;
      LAYER via ;
        RECT 541.750 499.160 542.010 499.420 ;
        RECT 542.900 497.800 543.160 498.060 ;
        RECT 540.600 471.620 540.860 471.880 ;
        RECT 542.440 471.620 542.700 471.880 ;
        RECT 540.600 80.620 540.860 80.880 ;
        RECT 1353.880 80.620 1354.140 80.880 ;
      LAYER met2 ;
        RECT 541.770 500.000 542.050 504.000 ;
        RECT 541.810 499.450 541.950 500.000 ;
        RECT 541.750 499.130 542.010 499.450 ;
        RECT 542.900 497.770 543.160 498.090 ;
        RECT 542.960 476.170 543.100 497.770 ;
        RECT 542.500 476.030 543.100 476.170 ;
        RECT 542.500 471.910 542.640 476.030 ;
        RECT 540.600 471.590 540.860 471.910 ;
        RECT 542.440 471.590 542.700 471.910 ;
        RECT 540.660 80.910 540.800 471.590 ;
        RECT 540.600 80.590 540.860 80.910 ;
        RECT 1353.880 80.590 1354.140 80.910 ;
        RECT 1353.940 1.770 1354.080 80.590 ;
        RECT 1356.030 1.770 1356.590 2.400 ;
        RECT 1353.940 1.630 1356.590 1.770 ;
        RECT 1356.030 -4.800 1356.590 1.630 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.150 500.000 543.430 504.000 ;
        RECT 543.190 498.850 543.330 500.000 ;
        RECT 543.190 498.710 543.560 498.850 ;
        RECT 543.420 491.485 543.560 498.710 ;
        RECT 543.350 491.115 543.630 491.485 ;
        RECT 1374.110 37.555 1374.390 37.925 ;
        RECT 1374.180 2.400 1374.320 37.555 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
      LAYER via2 ;
        RECT 543.350 491.160 543.630 491.440 ;
        RECT 1374.110 37.600 1374.390 37.880 ;
      LAYER met3 ;
        RECT 543.325 491.450 543.655 491.465 ;
        RECT 543.990 491.450 544.370 491.460 ;
        RECT 543.325 491.150 544.370 491.450 ;
        RECT 543.325 491.135 543.655 491.150 ;
        RECT 543.990 491.140 544.370 491.150 ;
        RECT 543.990 37.890 544.370 37.900 ;
        RECT 1374.085 37.890 1374.415 37.905 ;
        RECT 543.990 37.590 1374.415 37.890 ;
        RECT 543.990 37.580 544.370 37.590 ;
        RECT 1374.085 37.575 1374.415 37.590 ;
      LAYER via3 ;
        RECT 544.020 491.140 544.340 491.460 ;
        RECT 544.020 37.580 544.340 37.900 ;
      LAYER met4 ;
        RECT 544.015 491.135 544.345 491.465 ;
        RECT 544.030 37.905 544.330 491.135 ;
        RECT 544.015 37.575 544.345 37.905 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.530 500.000 544.810 504.000 ;
        RECT 544.570 499.645 544.710 500.000 ;
        RECT 544.500 499.275 544.780 499.645 ;
        RECT 1391.590 82.435 1391.870 82.805 ;
        RECT 1391.660 2.400 1391.800 82.435 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
      LAYER via2 ;
        RECT 544.500 499.320 544.780 499.600 ;
        RECT 1391.590 82.480 1391.870 82.760 ;
      LAYER met3 ;
        RECT 544.475 499.295 544.805 499.625 ;
        RECT 542.150 498.930 542.530 498.940 ;
        RECT 544.490 498.930 544.790 499.295 ;
        RECT 542.150 498.630 544.790 498.930 ;
        RECT 542.150 498.620 542.530 498.630 ;
        RECT 542.150 82.770 542.530 82.780 ;
        RECT 1391.565 82.770 1391.895 82.785 ;
        RECT 542.150 82.470 1391.895 82.770 ;
        RECT 542.150 82.460 542.530 82.470 ;
        RECT 1391.565 82.455 1391.895 82.470 ;
      LAYER via3 ;
        RECT 542.180 498.620 542.500 498.940 ;
        RECT 542.180 82.460 542.500 82.780 ;
      LAYER met4 ;
        RECT 542.175 498.615 542.505 498.945 ;
        RECT 542.190 82.785 542.490 498.615 ;
        RECT 542.175 82.455 542.505 82.785 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.860 499.700 546.180 499.760 ;
        RECT 545.030 499.560 546.180 499.700 ;
        RECT 545.030 496.640 545.170 499.560 ;
        RECT 545.860 499.500 546.180 499.560 ;
        RECT 1407.670 496.640 1407.990 496.700 ;
        RECT 545.030 496.500 1407.990 496.640 ;
        RECT 1407.670 496.440 1407.990 496.500 ;
      LAYER via ;
        RECT 545.890 499.500 546.150 499.760 ;
        RECT 1407.700 496.440 1407.960 496.700 ;
      LAYER met2 ;
        RECT 545.910 500.000 546.190 504.000 ;
        RECT 545.950 499.790 546.090 500.000 ;
        RECT 545.890 499.470 546.150 499.790 ;
        RECT 1407.700 496.410 1407.960 496.730 ;
        RECT 1407.760 1.770 1407.900 496.410 ;
        RECT 1409.390 1.770 1409.950 2.400 ;
        RECT 1407.760 1.630 1409.950 1.770 ;
        RECT 1409.390 -4.800 1409.950 1.630 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 547.010 498.480 547.330 498.740 ;
        RECT 547.100 498.060 547.240 498.480 ;
        RECT 547.010 497.800 547.330 498.060 ;
        RECT 546.550 89.660 546.870 89.720 ;
        RECT 1421.930 89.660 1422.250 89.720 ;
        RECT 546.550 89.520 1422.250 89.660 ;
        RECT 546.550 89.460 546.870 89.520 ;
        RECT 1421.930 89.460 1422.250 89.520 ;
      LAYER via ;
        RECT 547.040 498.480 547.300 498.740 ;
        RECT 547.040 497.800 547.300 498.060 ;
        RECT 546.580 89.460 546.840 89.720 ;
        RECT 1421.960 89.460 1422.220 89.720 ;
      LAYER met2 ;
        RECT 547.290 500.000 547.570 504.000 ;
        RECT 547.330 498.850 547.470 500.000 ;
        RECT 547.100 498.770 547.470 498.850 ;
        RECT 547.040 498.710 547.470 498.770 ;
        RECT 547.040 498.450 547.300 498.710 ;
        RECT 547.040 497.770 547.300 498.090 ;
        RECT 547.100 476.170 547.240 497.770 ;
        RECT 546.640 476.030 547.240 476.170 ;
        RECT 546.640 89.750 546.780 476.030 ;
        RECT 546.580 89.430 546.840 89.750 ;
        RECT 1421.960 89.430 1422.220 89.750 ;
        RECT 1422.020 82.870 1422.160 89.430 ;
        RECT 1422.020 82.730 1424.920 82.870 ;
        RECT 1424.780 1.770 1424.920 82.730 ;
        RECT 1426.870 1.770 1427.430 2.400 ;
        RECT 1424.780 1.630 1427.430 1.770 ;
        RECT 1426.870 -4.800 1427.430 1.630 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 548.620 500.860 548.940 501.120 ;
        RECT 547.470 498.000 547.790 498.060 ;
        RECT 548.710 498.000 548.850 500.860 ;
        RECT 547.470 497.860 548.850 498.000 ;
        RECT 547.470 497.800 547.790 497.860 ;
        RECT 546.090 489.840 546.410 489.900 ;
        RECT 547.470 489.840 547.790 489.900 ;
        RECT 546.090 489.700 547.790 489.840 ;
        RECT 546.090 489.640 546.410 489.700 ;
        RECT 547.470 489.640 547.790 489.700 ;
        RECT 545.630 89.320 545.950 89.380 ;
        RECT 1442.170 89.320 1442.490 89.380 ;
        RECT 545.630 89.180 1442.490 89.320 ;
        RECT 545.630 89.120 545.950 89.180 ;
        RECT 1442.170 89.120 1442.490 89.180 ;
      LAYER via ;
        RECT 548.650 500.860 548.910 501.120 ;
        RECT 547.500 497.800 547.760 498.060 ;
        RECT 546.120 489.640 546.380 489.900 ;
        RECT 547.500 489.640 547.760 489.900 ;
        RECT 545.660 89.120 545.920 89.380 ;
        RECT 1442.200 89.120 1442.460 89.380 ;
      LAYER met2 ;
        RECT 548.670 501.150 548.950 504.000 ;
        RECT 548.650 500.830 548.950 501.150 ;
        RECT 548.670 500.000 548.950 500.830 ;
        RECT 547.500 497.770 547.760 498.090 ;
        RECT 547.560 489.930 547.700 497.770 ;
        RECT 546.120 489.610 546.380 489.930 ;
        RECT 547.500 489.610 547.760 489.930 ;
        RECT 546.180 473.010 546.320 489.610 ;
        RECT 545.720 472.870 546.320 473.010 ;
        RECT 545.720 89.410 545.860 472.870 ;
        RECT 545.660 89.090 545.920 89.410 ;
        RECT 1442.200 89.090 1442.460 89.410 ;
        RECT 1442.260 82.870 1442.400 89.090 ;
        RECT 1442.260 82.730 1445.160 82.870 ;
        RECT 1445.020 2.400 1445.160 82.730 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 550.000 499.360 550.320 499.420 ;
        RECT 550.000 499.160 550.460 499.360 ;
        RECT 550.320 498.740 550.460 499.160 ;
        RECT 550.230 498.480 550.550 498.740 ;
        RECT 546.090 472.160 546.410 472.220 ;
        RECT 550.230 472.160 550.550 472.220 ;
        RECT 546.090 472.020 550.550 472.160 ;
        RECT 546.090 471.960 546.410 472.020 ;
        RECT 550.230 471.960 550.550 472.020 ;
        RECT 546.090 88.980 546.410 89.040 ;
        RECT 1462.870 88.980 1463.190 89.040 ;
        RECT 546.090 88.840 1463.190 88.980 ;
        RECT 546.090 88.780 546.410 88.840 ;
        RECT 1462.870 88.780 1463.190 88.840 ;
      LAYER via ;
        RECT 550.030 499.160 550.290 499.420 ;
        RECT 550.260 498.480 550.520 498.740 ;
        RECT 546.120 471.960 546.380 472.220 ;
        RECT 550.260 471.960 550.520 472.220 ;
        RECT 546.120 88.780 546.380 89.040 ;
        RECT 1462.900 88.780 1463.160 89.040 ;
      LAYER met2 ;
        RECT 550.050 500.000 550.330 504.000 ;
        RECT 550.090 499.450 550.230 500.000 ;
        RECT 550.030 499.130 550.290 499.450 ;
        RECT 550.260 498.450 550.520 498.770 ;
        RECT 550.320 472.250 550.460 498.450 ;
        RECT 546.120 471.930 546.380 472.250 ;
        RECT 550.260 471.930 550.520 472.250 ;
        RECT 546.180 89.070 546.320 471.930 ;
        RECT 546.120 88.750 546.380 89.070 ;
        RECT 1462.900 88.750 1463.160 89.070 ;
        RECT 1462.960 2.400 1463.100 88.750 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.430 500.000 551.710 504.000 ;
        RECT 551.470 499.815 551.610 500.000 ;
        RECT 551.400 499.445 551.680 499.815 ;
        RECT 1476.690 86.515 1476.970 86.885 ;
        RECT 1476.760 82.870 1476.900 86.515 ;
        RECT 1476.760 82.730 1478.280 82.870 ;
        RECT 1478.140 1.770 1478.280 82.730 ;
        RECT 1480.230 1.770 1480.790 2.400 ;
        RECT 1478.140 1.630 1480.790 1.770 ;
        RECT 1480.230 -4.800 1480.790 1.630 ;
      LAYER via2 ;
        RECT 551.400 499.490 551.680 499.770 ;
        RECT 1476.690 86.560 1476.970 86.840 ;
      LAYER met3 ;
        RECT 547.670 500.290 548.050 500.300 ;
        RECT 550.700 500.290 551.690 500.460 ;
        RECT 547.670 500.160 551.690 500.290 ;
        RECT 547.670 499.990 551.000 500.160 ;
        RECT 547.670 499.980 548.050 499.990 ;
        RECT 551.390 499.795 551.690 500.160 ;
        RECT 551.375 499.465 551.705 499.795 ;
        RECT 547.670 86.850 548.050 86.860 ;
        RECT 1476.665 86.850 1476.995 86.865 ;
        RECT 547.670 86.550 1476.995 86.850 ;
        RECT 547.670 86.540 548.050 86.550 ;
        RECT 1476.665 86.535 1476.995 86.550 ;
      LAYER via3 ;
        RECT 547.700 499.980 548.020 500.300 ;
        RECT 547.700 86.540 548.020 86.860 ;
      LAYER met4 ;
        RECT 547.695 499.975 548.025 500.305 ;
        RECT 547.710 86.865 548.010 499.975 ;
        RECT 547.695 86.535 548.025 86.865 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.760 499.500 553.080 499.760 ;
        RECT 552.850 499.080 552.990 499.500 ;
        RECT 552.850 498.880 553.310 499.080 ;
        RECT 552.990 498.820 553.310 498.880 ;
        RECT 552.990 496.300 553.310 496.360 ;
        RECT 1497.370 496.300 1497.690 496.360 ;
        RECT 552.990 496.160 1497.690 496.300 ;
        RECT 552.990 496.100 553.310 496.160 ;
        RECT 1497.370 496.100 1497.690 496.160 ;
      LAYER via ;
        RECT 552.790 499.500 553.050 499.760 ;
        RECT 553.020 498.820 553.280 499.080 ;
        RECT 553.020 496.100 553.280 496.360 ;
        RECT 1497.400 496.100 1497.660 496.360 ;
      LAYER met2 ;
        RECT 552.810 500.000 553.090 504.000 ;
        RECT 552.850 499.790 552.990 500.000 ;
        RECT 552.790 499.470 553.050 499.790 ;
        RECT 553.020 498.790 553.280 499.110 ;
        RECT 553.080 496.390 553.220 498.790 ;
        RECT 553.020 496.070 553.280 496.390 ;
        RECT 1497.400 496.070 1497.660 496.390 ;
        RECT 1497.460 17.410 1497.600 496.070 ;
        RECT 1497.460 17.270 1498.520 17.410 ;
        RECT 1498.380 2.400 1498.520 17.270 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.660 500.380 490.980 500.440 ;
        RECT 489.830 500.240 490.980 500.380 ;
        RECT 489.830 497.720 489.970 500.240 ;
        RECT 490.660 500.180 490.980 500.240 ;
        RECT 489.830 497.520 490.290 497.720 ;
        RECT 489.970 497.460 490.290 497.520 ;
        RECT 489.970 47.500 490.290 47.560 ;
        RECT 700.190 47.500 700.510 47.560 ;
        RECT 489.970 47.360 700.510 47.500 ;
        RECT 489.970 47.300 490.290 47.360 ;
        RECT 700.190 47.300 700.510 47.360 ;
      LAYER via ;
        RECT 490.690 500.180 490.950 500.440 ;
        RECT 490.000 497.460 490.260 497.720 ;
        RECT 490.000 47.300 490.260 47.560 ;
        RECT 700.220 47.300 700.480 47.560 ;
      LAYER met2 ;
        RECT 490.710 500.470 490.990 504.000 ;
        RECT 490.690 500.150 490.990 500.470 ;
        RECT 490.710 500.000 490.990 500.150 ;
        RECT 490.000 497.430 490.260 497.750 ;
        RECT 490.060 47.590 490.200 497.430 ;
        RECT 490.000 47.270 490.260 47.590 ;
        RECT 700.220 47.270 700.480 47.590 ;
        RECT 700.280 2.400 700.420 47.270 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 553.450 95.440 553.770 95.500 ;
        RECT 1511.170 95.440 1511.490 95.500 ;
        RECT 553.450 95.300 1511.490 95.440 ;
        RECT 553.450 95.240 553.770 95.300 ;
        RECT 1511.170 95.240 1511.490 95.300 ;
      LAYER via ;
        RECT 553.480 95.240 553.740 95.500 ;
        RECT 1511.200 95.240 1511.460 95.500 ;
      LAYER met2 ;
        RECT 554.190 500.000 554.470 504.000 ;
        RECT 554.230 499.815 554.370 500.000 ;
        RECT 554.160 499.445 554.440 499.815 ;
        RECT 553.930 498.595 554.210 498.965 ;
        RECT 554.000 490.860 554.140 498.595 ;
        RECT 553.540 490.720 554.140 490.860 ;
        RECT 553.540 95.530 553.680 490.720 ;
        RECT 553.480 95.210 553.740 95.530 ;
        RECT 1511.200 95.210 1511.460 95.530 ;
        RECT 1511.260 82.870 1511.400 95.210 ;
        RECT 1511.260 82.730 1516.000 82.870 ;
        RECT 1515.860 2.400 1516.000 82.730 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
      LAYER via2 ;
        RECT 554.160 499.490 554.440 499.770 ;
        RECT 553.930 498.640 554.210 498.920 ;
      LAYER met3 ;
        RECT 554.135 499.465 554.465 499.795 ;
        RECT 554.150 498.945 554.450 499.465 ;
        RECT 553.905 498.630 554.450 498.945 ;
        RECT 553.905 498.615 554.235 498.630 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 555.520 499.500 555.840 499.760 ;
        RECT 555.610 498.400 555.750 499.500 ;
        RECT 555.610 498.200 556.070 498.400 ;
        RECT 555.750 498.140 556.070 498.200 ;
        RECT 553.910 490.180 554.230 490.240 ;
        RECT 555.750 490.180 556.070 490.240 ;
        RECT 553.910 490.040 556.070 490.180 ;
        RECT 553.910 489.980 554.230 490.040 ;
        RECT 555.750 489.980 556.070 490.040 ;
        RECT 553.910 95.100 554.230 95.160 ;
        RECT 1531.870 95.100 1532.190 95.160 ;
        RECT 553.910 94.960 1532.190 95.100 ;
        RECT 553.910 94.900 554.230 94.960 ;
        RECT 1531.870 94.900 1532.190 94.960 ;
      LAYER via ;
        RECT 555.550 499.500 555.810 499.760 ;
        RECT 555.780 498.140 556.040 498.400 ;
        RECT 553.940 489.980 554.200 490.240 ;
        RECT 555.780 489.980 556.040 490.240 ;
        RECT 553.940 94.900 554.200 95.160 ;
        RECT 1531.900 94.900 1532.160 95.160 ;
      LAYER met2 ;
        RECT 555.570 500.000 555.850 504.000 ;
        RECT 555.610 499.790 555.750 500.000 ;
        RECT 555.550 499.470 555.810 499.790 ;
        RECT 555.780 498.110 556.040 498.430 ;
        RECT 555.840 490.270 555.980 498.110 ;
        RECT 553.940 489.950 554.200 490.270 ;
        RECT 555.780 489.950 556.040 490.270 ;
        RECT 554.000 95.190 554.140 489.950 ;
        RECT 553.940 94.870 554.200 95.190 ;
        RECT 1531.900 94.870 1532.160 95.190 ;
        RECT 1531.960 1.770 1532.100 94.870 ;
        RECT 1533.590 1.770 1534.150 2.400 ;
        RECT 1531.960 1.630 1534.150 1.770 ;
        RECT 1533.590 -4.800 1534.150 1.630 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.950 500.000 557.230 504.000 ;
        RECT 556.990 498.680 557.130 500.000 ;
        RECT 556.990 498.540 557.360 498.680 ;
        RECT 557.220 491.485 557.360 498.540 ;
        RECT 557.150 491.115 557.430 491.485 ;
        RECT 1551.210 32.115 1551.490 32.485 ;
        RECT 1551.280 2.400 1551.420 32.115 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
      LAYER via2 ;
        RECT 557.150 491.160 557.430 491.440 ;
        RECT 1551.210 32.160 1551.490 32.440 ;
      LAYER met3 ;
        RECT 557.125 491.460 557.455 491.465 ;
        RECT 556.870 491.450 557.455 491.460 ;
        RECT 556.670 491.150 557.455 491.450 ;
        RECT 556.870 491.140 557.455 491.150 ;
        RECT 557.125 491.135 557.455 491.140 ;
        RECT 556.870 32.450 557.250 32.460 ;
        RECT 1551.185 32.450 1551.515 32.465 ;
        RECT 556.870 32.150 1551.515 32.450 ;
        RECT 556.870 32.140 557.250 32.150 ;
        RECT 1551.185 32.135 1551.515 32.150 ;
      LAYER via3 ;
        RECT 556.900 491.140 557.220 491.460 ;
        RECT 556.900 32.140 557.220 32.460 ;
      LAYER met4 ;
        RECT 556.895 491.135 557.225 491.465 ;
        RECT 556.910 32.465 557.210 491.135 ;
        RECT 556.895 32.135 557.225 32.465 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.330 500.000 558.610 504.000 ;
        RECT 558.370 499.645 558.510 500.000 ;
        RECT 558.300 499.275 558.580 499.645 ;
        RECT 1569.150 31.435 1569.430 31.805 ;
        RECT 1569.220 2.400 1569.360 31.435 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
      LAYER via2 ;
        RECT 558.300 499.320 558.580 499.600 ;
        RECT 1569.150 31.480 1569.430 31.760 ;
      LAYER met3 ;
        RECT 558.275 499.610 558.605 499.625 ;
        RECT 558.275 499.295 558.820 499.610 ;
        RECT 557.790 498.930 558.170 498.940 ;
        RECT 558.520 498.930 558.820 499.295 ;
        RECT 557.790 498.630 558.820 498.930 ;
        RECT 557.790 498.620 558.170 498.630 ;
        RECT 557.790 31.770 558.170 31.780 ;
        RECT 1569.125 31.770 1569.455 31.785 ;
        RECT 557.790 31.470 1569.455 31.770 ;
        RECT 557.790 31.460 558.170 31.470 ;
        RECT 1569.125 31.455 1569.455 31.470 ;
      LAYER via3 ;
        RECT 557.820 498.620 558.140 498.940 ;
        RECT 557.820 31.460 558.140 31.780 ;
      LAYER met4 ;
        RECT 557.815 498.615 558.145 498.945 ;
        RECT 557.830 31.785 558.130 498.615 ;
        RECT 557.815 31.455 558.145 31.785 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.660 499.500 559.980 499.760 ;
        RECT 559.750 499.360 559.890 499.500 ;
        RECT 559.750 499.220 560.120 499.360 ;
        RECT 559.980 498.740 560.120 499.220 ;
        RECT 559.890 498.480 560.210 498.740 ;
        RECT 559.890 495.960 560.210 496.020 ;
        RECT 1580.170 495.960 1580.490 496.020 ;
        RECT 559.890 495.820 1580.490 495.960 ;
        RECT 559.890 495.760 560.210 495.820 ;
        RECT 1580.170 495.760 1580.490 495.820 ;
        RECT 1580.170 16.900 1580.490 16.960 ;
        RECT 1586.610 16.900 1586.930 16.960 ;
        RECT 1580.170 16.760 1586.930 16.900 ;
        RECT 1580.170 16.700 1580.490 16.760 ;
        RECT 1586.610 16.700 1586.930 16.760 ;
      LAYER via ;
        RECT 559.690 499.500 559.950 499.760 ;
        RECT 559.920 498.480 560.180 498.740 ;
        RECT 559.920 495.760 560.180 496.020 ;
        RECT 1580.200 495.760 1580.460 496.020 ;
        RECT 1580.200 16.700 1580.460 16.960 ;
        RECT 1586.640 16.700 1586.900 16.960 ;
      LAYER met2 ;
        RECT 559.710 500.000 559.990 504.000 ;
        RECT 559.750 499.790 559.890 500.000 ;
        RECT 559.690 499.470 559.950 499.790 ;
        RECT 559.920 498.450 560.180 498.770 ;
        RECT 559.980 496.050 560.120 498.450 ;
        RECT 559.920 495.730 560.180 496.050 ;
        RECT 1580.200 495.730 1580.460 496.050 ;
        RECT 1580.260 16.990 1580.400 495.730 ;
        RECT 1580.200 16.670 1580.460 16.990 ;
        RECT 1586.640 16.670 1586.900 16.990 ;
        RECT 1586.700 2.400 1586.840 16.670 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 561.040 499.160 561.360 499.420 ;
        RECT 561.130 498.740 561.270 499.160 ;
        RECT 561.130 498.540 561.590 498.740 ;
        RECT 561.270 498.480 561.590 498.540 ;
        RECT 559.890 491.880 560.210 491.940 ;
        RECT 561.270 491.880 561.590 491.940 ;
        RECT 559.890 491.740 561.590 491.880 ;
        RECT 559.890 491.680 560.210 491.740 ;
        RECT 561.270 491.680 561.590 491.740 ;
        RECT 559.890 94.760 560.210 94.820 ;
        RECT 1600.870 94.760 1601.190 94.820 ;
        RECT 559.890 94.620 1601.190 94.760 ;
        RECT 559.890 94.560 560.210 94.620 ;
        RECT 1600.870 94.560 1601.190 94.620 ;
      LAYER via ;
        RECT 561.070 499.160 561.330 499.420 ;
        RECT 561.300 498.480 561.560 498.740 ;
        RECT 559.920 491.680 560.180 491.940 ;
        RECT 561.300 491.680 561.560 491.940 ;
        RECT 559.920 94.560 560.180 94.820 ;
        RECT 1600.900 94.560 1601.160 94.820 ;
      LAYER met2 ;
        RECT 561.090 500.000 561.370 504.000 ;
        RECT 561.130 499.450 561.270 500.000 ;
        RECT 561.070 499.130 561.330 499.450 ;
        RECT 561.300 498.450 561.560 498.770 ;
        RECT 561.360 491.970 561.500 498.450 ;
        RECT 559.920 491.650 560.180 491.970 ;
        RECT 561.300 491.650 561.560 491.970 ;
        RECT 559.980 94.850 560.120 491.650 ;
        RECT 559.920 94.530 560.180 94.850 ;
        RECT 1600.900 94.530 1601.160 94.850 ;
        RECT 1600.960 82.870 1601.100 94.530 ;
        RECT 1600.960 82.730 1602.480 82.870 ;
        RECT 1602.340 1.770 1602.480 82.730 ;
        RECT 1604.430 1.770 1604.990 2.400 ;
        RECT 1602.340 1.630 1604.990 1.770 ;
        RECT 1604.430 -4.800 1604.990 1.630 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 561.270 491.200 561.590 491.260 ;
        RECT 562.650 491.200 562.970 491.260 ;
        RECT 561.270 491.060 562.970 491.200 ;
        RECT 561.270 491.000 561.590 491.060 ;
        RECT 562.650 491.000 562.970 491.060 ;
        RECT 558.970 471.480 559.290 471.540 ;
        RECT 561.730 471.480 562.050 471.540 ;
        RECT 558.970 471.340 562.050 471.480 ;
        RECT 558.970 471.280 559.290 471.340 ;
        RECT 561.730 471.280 562.050 471.340 ;
        RECT 558.970 45.800 559.290 45.860 ;
        RECT 1622.030 45.800 1622.350 45.860 ;
        RECT 558.970 45.660 1622.350 45.800 ;
        RECT 558.970 45.600 559.290 45.660 ;
        RECT 1622.030 45.600 1622.350 45.660 ;
      LAYER via ;
        RECT 561.300 491.000 561.560 491.260 ;
        RECT 562.680 491.000 562.940 491.260 ;
        RECT 559.000 471.280 559.260 471.540 ;
        RECT 561.760 471.280 562.020 471.540 ;
        RECT 559.000 45.600 559.260 45.860 ;
        RECT 1622.060 45.600 1622.320 45.860 ;
      LAYER met2 ;
        RECT 562.470 500.000 562.750 504.000 ;
        RECT 562.510 499.475 562.650 500.000 ;
        RECT 562.440 499.105 562.720 499.475 ;
        RECT 562.670 497.235 562.950 497.605 ;
        RECT 562.740 491.290 562.880 497.235 ;
        RECT 561.300 490.970 561.560 491.290 ;
        RECT 562.680 490.970 562.940 491.290 ;
        RECT 561.360 473.690 561.500 490.970 ;
        RECT 561.360 473.550 561.960 473.690 ;
        RECT 561.820 471.570 561.960 473.550 ;
        RECT 559.000 471.250 559.260 471.570 ;
        RECT 561.760 471.250 562.020 471.570 ;
        RECT 559.060 45.890 559.200 471.250 ;
        RECT 559.000 45.570 559.260 45.890 ;
        RECT 1622.060 45.570 1622.320 45.890 ;
        RECT 1622.120 2.400 1622.260 45.570 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
      LAYER via2 ;
        RECT 562.440 499.150 562.720 499.430 ;
        RECT 562.670 497.280 562.950 497.560 ;
      LAYER met3 ;
        RECT 562.415 499.125 562.745 499.455 ;
        RECT 562.430 497.585 562.730 499.125 ;
        RECT 562.430 497.270 562.975 497.585 ;
        RECT 562.645 497.255 562.975 497.270 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 563.800 499.500 564.120 499.760 ;
        RECT 563.890 498.740 564.030 499.500 ;
        RECT 563.890 498.540 564.350 498.740 ;
        RECT 564.030 498.480 564.350 498.540 ;
      LAYER via ;
        RECT 563.830 499.500 564.090 499.760 ;
        RECT 564.060 498.480 564.320 498.740 ;
      LAYER met2 ;
        RECT 563.850 500.000 564.130 504.000 ;
        RECT 563.890 499.790 564.030 500.000 ;
        RECT 563.830 499.470 564.090 499.790 ;
        RECT 564.060 498.450 564.320 498.770 ;
        RECT 564.120 492.165 564.260 498.450 ;
        RECT 564.050 491.795 564.330 492.165 ;
        RECT 1639.990 51.835 1640.270 52.205 ;
        RECT 1640.060 2.400 1640.200 51.835 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
      LAYER via2 ;
        RECT 564.050 491.840 564.330 492.120 ;
        RECT 1639.990 51.880 1640.270 52.160 ;
      LAYER met3 ;
        RECT 564.025 492.130 564.355 492.145 ;
        RECT 565.150 492.130 565.530 492.140 ;
        RECT 564.025 491.830 565.530 492.130 ;
        RECT 564.025 491.815 564.355 491.830 ;
        RECT 565.150 491.820 565.530 491.830 ;
        RECT 565.150 52.170 565.530 52.180 ;
        RECT 1639.965 52.170 1640.295 52.185 ;
        RECT 565.150 51.870 1640.295 52.170 ;
        RECT 565.150 51.860 565.530 51.870 ;
        RECT 1639.965 51.855 1640.295 51.870 ;
      LAYER via3 ;
        RECT 565.180 491.820 565.500 492.140 ;
        RECT 565.180 51.860 565.500 52.180 ;
      LAYER met4 ;
        RECT 565.175 491.815 565.505 492.145 ;
        RECT 565.190 52.185 565.490 491.815 ;
        RECT 565.175 51.855 565.505 52.185 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.230 500.000 565.510 504.000 ;
        RECT 565.270 499.815 565.410 500.000 ;
        RECT 565.200 499.445 565.480 499.815 ;
        RECT 1656.090 94.675 1656.370 95.045 ;
        RECT 1656.160 1.770 1656.300 94.675 ;
        RECT 1657.790 1.770 1658.350 2.400 ;
        RECT 1656.160 1.630 1658.350 1.770 ;
        RECT 1657.790 -4.800 1658.350 1.630 ;
      LAYER via2 ;
        RECT 565.200 499.490 565.480 499.770 ;
        RECT 1656.090 94.720 1656.370 95.000 ;
      LAYER met3 ;
        RECT 565.175 499.465 565.505 499.795 ;
        RECT 563.310 498.930 563.690 498.940 ;
        RECT 565.190 498.930 565.490 499.465 ;
        RECT 563.310 498.630 565.490 498.930 ;
        RECT 563.310 498.620 563.690 498.630 ;
        RECT 563.310 95.010 563.690 95.020 ;
        RECT 1656.065 95.010 1656.395 95.025 ;
        RECT 563.310 94.710 1656.395 95.010 ;
        RECT 563.310 94.700 563.690 94.710 ;
        RECT 1656.065 94.695 1656.395 94.710 ;
      LAYER via3 ;
        RECT 563.340 498.620 563.660 498.940 ;
        RECT 563.340 94.700 563.660 95.020 ;
      LAYER met4 ;
        RECT 563.335 498.615 563.665 498.945 ;
        RECT 563.350 95.025 563.650 498.615 ;
        RECT 563.335 94.695 563.665 95.025 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.560 498.820 566.880 499.080 ;
        RECT 566.650 498.340 566.790 498.820 ;
        RECT 567.250 498.340 567.570 498.400 ;
        RECT 566.650 498.200 567.570 498.340 ;
        RECT 567.250 498.140 567.570 498.200 ;
        RECT 618.770 495.620 619.090 495.680 ;
        RECT 1669.870 495.620 1670.190 495.680 ;
        RECT 618.770 495.480 1670.190 495.620 ;
        RECT 618.770 495.420 619.090 495.480 ;
        RECT 1669.870 495.420 1670.190 495.480 ;
        RECT 567.250 493.240 567.570 493.300 ;
        RECT 618.770 493.240 619.090 493.300 ;
        RECT 567.250 493.100 619.090 493.240 ;
        RECT 567.250 493.040 567.570 493.100 ;
        RECT 618.770 493.040 619.090 493.100 ;
      LAYER via ;
        RECT 566.590 498.820 566.850 499.080 ;
        RECT 567.280 498.140 567.540 498.400 ;
        RECT 618.800 495.420 619.060 495.680 ;
        RECT 1669.900 495.420 1670.160 495.680 ;
        RECT 567.280 493.040 567.540 493.300 ;
        RECT 618.800 493.040 619.060 493.300 ;
      LAYER met2 ;
        RECT 566.610 500.000 566.890 504.000 ;
        RECT 566.650 499.110 566.790 500.000 ;
        RECT 566.590 498.790 566.850 499.110 ;
        RECT 567.280 498.110 567.540 498.430 ;
        RECT 567.340 493.330 567.480 498.110 ;
        RECT 618.800 495.390 619.060 495.710 ;
        RECT 1669.900 495.390 1670.160 495.710 ;
        RECT 618.860 493.330 619.000 495.390 ;
        RECT 567.280 493.010 567.540 493.330 ;
        RECT 618.800 493.010 619.060 493.330 ;
        RECT 1669.960 82.870 1670.100 495.390 ;
        RECT 1669.960 82.730 1673.320 82.870 ;
        RECT 1673.180 1.770 1673.320 82.730 ;
        RECT 1675.270 1.770 1675.830 2.400 ;
        RECT 1673.180 1.630 1675.830 1.770 ;
        RECT 1675.270 -4.800 1675.830 1.630 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 492.040 499.360 492.360 499.420 ;
        RECT 491.900 499.160 492.360 499.360 ;
        RECT 491.900 498.740 492.040 499.160 ;
        RECT 491.810 498.480 492.130 498.740 ;
        RECT 491.810 102.580 492.130 102.640 ;
        RECT 718.130 102.580 718.450 102.640 ;
        RECT 491.810 102.440 718.450 102.580 ;
        RECT 491.810 102.380 492.130 102.440 ;
        RECT 718.130 102.380 718.450 102.440 ;
      LAYER via ;
        RECT 492.070 499.160 492.330 499.420 ;
        RECT 491.840 498.480 492.100 498.740 ;
        RECT 491.840 102.380 492.100 102.640 ;
        RECT 718.160 102.380 718.420 102.640 ;
      LAYER met2 ;
        RECT 492.090 500.000 492.370 504.000 ;
        RECT 492.130 499.450 492.270 500.000 ;
        RECT 492.070 499.130 492.330 499.450 ;
        RECT 491.840 498.450 492.100 498.770 ;
        RECT 491.900 102.670 492.040 498.450 ;
        RECT 491.840 102.350 492.100 102.670 ;
        RECT 718.160 102.350 718.420 102.670 ;
        RECT 718.220 34.570 718.360 102.350 ;
        RECT 717.760 34.430 718.360 34.570 ;
        RECT 717.760 2.400 717.900 34.430 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 567.940 499.160 568.260 499.420 ;
        RECT 568.030 498.740 568.170 499.160 ;
        RECT 567.710 498.540 568.170 498.740 ;
        RECT 567.710 498.480 568.030 498.540 ;
        RECT 567.710 101.900 568.030 101.960 ;
        RECT 1690.570 101.900 1690.890 101.960 ;
        RECT 567.710 101.760 1690.890 101.900 ;
        RECT 567.710 101.700 568.030 101.760 ;
        RECT 1690.570 101.700 1690.890 101.760 ;
      LAYER via ;
        RECT 567.970 499.160 568.230 499.420 ;
        RECT 567.740 498.480 568.000 498.740 ;
        RECT 567.740 101.700 568.000 101.960 ;
        RECT 1690.600 101.700 1690.860 101.960 ;
      LAYER met2 ;
        RECT 567.990 500.000 568.270 504.000 ;
        RECT 568.030 499.450 568.170 500.000 ;
        RECT 567.970 499.130 568.230 499.450 ;
        RECT 567.740 498.450 568.000 498.770 ;
        RECT 567.800 101.990 567.940 498.450 ;
        RECT 567.740 101.670 568.000 101.990 ;
        RECT 1690.600 101.670 1690.860 101.990 ;
        RECT 1690.660 82.870 1690.800 101.670 ;
        RECT 1690.660 82.730 1693.560 82.870 ;
        RECT 1693.420 2.400 1693.560 82.730 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 569.320 499.500 569.640 499.760 ;
        RECT 569.410 499.020 569.550 499.500 ;
        RECT 569.410 498.880 569.780 499.020 ;
        RECT 565.870 496.980 566.190 497.040 ;
        RECT 569.640 496.980 569.780 498.880 ;
        RECT 565.870 496.840 569.780 496.980 ;
        RECT 565.870 496.780 566.190 496.840 ;
        RECT 565.870 51.580 566.190 51.640 ;
        RECT 1704.830 51.580 1705.150 51.640 ;
        RECT 565.870 51.440 1705.150 51.580 ;
        RECT 565.870 51.380 566.190 51.440 ;
        RECT 1704.830 51.380 1705.150 51.440 ;
        RECT 1704.830 16.900 1705.150 16.960 ;
        RECT 1710.810 16.900 1711.130 16.960 ;
        RECT 1704.830 16.760 1711.130 16.900 ;
        RECT 1704.830 16.700 1705.150 16.760 ;
        RECT 1710.810 16.700 1711.130 16.760 ;
      LAYER via ;
        RECT 569.350 499.500 569.610 499.760 ;
        RECT 565.900 496.780 566.160 497.040 ;
        RECT 565.900 51.380 566.160 51.640 ;
        RECT 1704.860 51.380 1705.120 51.640 ;
        RECT 1704.860 16.700 1705.120 16.960 ;
        RECT 1710.840 16.700 1711.100 16.960 ;
      LAYER met2 ;
        RECT 569.370 500.000 569.650 504.000 ;
        RECT 569.410 499.790 569.550 500.000 ;
        RECT 569.350 499.470 569.610 499.790 ;
        RECT 565.900 496.750 566.160 497.070 ;
        RECT 565.960 51.670 566.100 496.750 ;
        RECT 565.900 51.350 566.160 51.670 ;
        RECT 1704.860 51.350 1705.120 51.670 ;
        RECT 1704.920 16.990 1705.060 51.350 ;
        RECT 1704.860 16.670 1705.120 16.990 ;
        RECT 1710.840 16.670 1711.100 16.990 ;
        RECT 1710.900 2.400 1711.040 16.670 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.750 500.000 571.030 504.000 ;
        RECT 570.790 499.645 570.930 500.000 ;
        RECT 570.720 499.275 571.000 499.645 ;
        RECT 1726.470 51.155 1726.750 51.525 ;
        RECT 1726.540 1.770 1726.680 51.155 ;
        RECT 1728.630 1.770 1729.190 2.400 ;
        RECT 1726.540 1.630 1729.190 1.770 ;
        RECT 1728.630 -4.800 1729.190 1.630 ;
      LAYER via2 ;
        RECT 570.720 499.320 571.000 499.600 ;
        RECT 1726.470 51.200 1726.750 51.480 ;
      LAYER met3 ;
        RECT 570.695 499.620 571.025 499.625 ;
        RECT 570.670 499.610 571.050 499.620 ;
        RECT 570.670 499.310 571.480 499.610 ;
        RECT 570.670 499.300 571.050 499.310 ;
        RECT 570.695 499.295 571.025 499.300 ;
        RECT 570.670 51.490 571.050 51.500 ;
        RECT 1726.445 51.490 1726.775 51.505 ;
        RECT 570.670 51.190 1726.775 51.490 ;
        RECT 570.670 51.180 571.050 51.190 ;
        RECT 1726.445 51.175 1726.775 51.190 ;
      LAYER via3 ;
        RECT 570.700 499.300 571.020 499.620 ;
        RECT 570.700 51.180 571.020 51.500 ;
      LAYER met4 ;
        RECT 570.695 499.295 571.025 499.625 ;
        RECT 570.710 51.505 571.010 499.295 ;
        RECT 570.695 51.175 571.025 51.505 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.130 500.000 572.410 504.000 ;
        RECT 572.170 499.815 572.310 500.000 ;
        RECT 572.100 499.445 572.380 499.815 ;
        RECT 1746.250 57.955 1746.530 58.325 ;
        RECT 1746.320 2.400 1746.460 57.955 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
      LAYER via2 ;
        RECT 572.100 499.490 572.380 499.770 ;
        RECT 1746.250 58.000 1746.530 58.280 ;
      LAYER met3 ;
        RECT 572.075 499.465 572.405 499.795 ;
        RECT 569.750 498.930 570.130 498.940 ;
        RECT 572.090 498.930 572.390 499.465 ;
        RECT 569.750 498.630 572.390 498.930 ;
        RECT 569.750 498.620 570.130 498.630 ;
        RECT 569.750 58.290 570.130 58.300 ;
        RECT 1746.225 58.290 1746.555 58.305 ;
        RECT 569.750 57.990 1746.555 58.290 ;
        RECT 569.750 57.980 570.130 57.990 ;
        RECT 1746.225 57.975 1746.555 57.990 ;
      LAYER via3 ;
        RECT 569.780 498.620 570.100 498.940 ;
        RECT 569.780 57.980 570.100 58.300 ;
      LAYER met4 ;
        RECT 569.775 498.615 570.105 498.945 ;
        RECT 569.790 58.305 570.090 498.615 ;
        RECT 569.775 57.975 570.105 58.305 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.610 495.620 574.930 495.680 ;
        RECT 574.610 495.480 617.620 495.620 ;
        RECT 574.610 495.420 574.930 495.480 ;
        RECT 617.480 495.280 617.620 495.480 ;
        RECT 1759.570 495.280 1759.890 495.340 ;
        RECT 617.480 495.140 1759.890 495.280 ;
        RECT 1759.570 495.080 1759.890 495.140 ;
      LAYER via ;
        RECT 574.640 495.420 574.900 495.680 ;
        RECT 1759.600 495.080 1759.860 495.340 ;
      LAYER met2 ;
        RECT 573.510 500.000 573.790 504.000 ;
        RECT 573.550 498.965 573.690 500.000 ;
        RECT 573.480 498.595 573.760 498.965 ;
        RECT 574.630 497.915 574.910 498.285 ;
        RECT 574.700 495.710 574.840 497.915 ;
        RECT 574.640 495.390 574.900 495.710 ;
        RECT 1759.600 495.050 1759.860 495.370 ;
        RECT 1759.660 82.870 1759.800 495.050 ;
        RECT 1759.660 82.730 1764.400 82.870 ;
        RECT 1764.260 2.400 1764.400 82.730 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
      LAYER via2 ;
        RECT 573.480 498.640 573.760 498.920 ;
        RECT 574.630 497.960 574.910 498.240 ;
      LAYER met3 ;
        RECT 573.455 498.615 573.785 498.945 ;
        RECT 573.470 498.250 573.770 498.615 ;
        RECT 574.605 498.250 574.935 498.265 ;
        RECT 573.470 497.950 574.935 498.250 ;
        RECT 574.605 497.935 574.935 497.950 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.840 499.160 575.160 499.420 ;
        RECT 573.690 498.340 574.010 498.400 ;
        RECT 574.930 498.340 575.070 499.160 ;
        RECT 573.690 498.200 575.070 498.340 ;
        RECT 573.690 498.140 574.010 498.200 ;
        RECT 573.690 101.560 574.010 101.620 ;
        RECT 1780.270 101.560 1780.590 101.620 ;
        RECT 573.690 101.420 1780.590 101.560 ;
        RECT 573.690 101.360 574.010 101.420 ;
        RECT 1780.270 101.360 1780.590 101.420 ;
      LAYER via ;
        RECT 574.870 499.160 575.130 499.420 ;
        RECT 573.720 498.140 573.980 498.400 ;
        RECT 573.720 101.360 573.980 101.620 ;
        RECT 1780.300 101.360 1780.560 101.620 ;
      LAYER met2 ;
        RECT 574.890 500.000 575.170 504.000 ;
        RECT 574.930 499.450 575.070 500.000 ;
        RECT 574.870 499.130 575.130 499.450 ;
        RECT 573.720 498.110 573.980 498.430 ;
        RECT 573.780 101.650 573.920 498.110 ;
        RECT 573.720 101.330 573.980 101.650 ;
        RECT 1780.300 101.330 1780.560 101.650 ;
        RECT 1780.360 82.870 1780.500 101.330 ;
        RECT 1780.360 82.730 1781.880 82.870 ;
        RECT 1781.740 2.400 1781.880 82.730 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 572.770 471.820 573.090 471.880 ;
        RECT 576.910 471.820 577.230 471.880 ;
        RECT 572.770 471.680 577.230 471.820 ;
        RECT 572.770 471.620 573.090 471.680 ;
        RECT 576.910 471.620 577.230 471.680 ;
        RECT 572.770 58.720 573.090 58.780 ;
        RECT 1797.290 58.720 1797.610 58.780 ;
        RECT 572.770 58.580 1797.610 58.720 ;
        RECT 572.770 58.520 573.090 58.580 ;
        RECT 1797.290 58.520 1797.610 58.580 ;
      LAYER via ;
        RECT 572.800 471.620 573.060 471.880 ;
        RECT 576.940 471.620 577.200 471.880 ;
        RECT 572.800 58.520 573.060 58.780 ;
        RECT 1797.320 58.520 1797.580 58.780 ;
      LAYER met2 ;
        RECT 576.270 500.000 576.550 504.000 ;
        RECT 576.310 498.850 576.450 500.000 ;
        RECT 576.310 498.710 576.680 498.850 ;
        RECT 576.540 473.690 576.680 498.710 ;
        RECT 576.540 473.550 577.140 473.690 ;
        RECT 577.000 471.910 577.140 473.550 ;
        RECT 572.800 471.590 573.060 471.910 ;
        RECT 576.940 471.590 577.200 471.910 ;
        RECT 572.860 58.810 573.000 471.590 ;
        RECT 572.800 58.490 573.060 58.810 ;
        RECT 1797.320 58.490 1797.580 58.810 ;
        RECT 1797.380 1.770 1797.520 58.490 ;
        RECT 1799.470 1.770 1800.030 2.400 ;
        RECT 1797.380 1.630 1800.030 1.770 ;
        RECT 1799.470 -4.800 1800.030 1.630 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.150 472.160 574.470 472.220 ;
        RECT 577.370 472.160 577.690 472.220 ;
        RECT 574.150 472.020 577.690 472.160 ;
        RECT 574.150 471.960 574.470 472.020 ;
        RECT 577.370 471.960 577.690 472.020 ;
        RECT 574.150 101.220 574.470 101.280 ;
        RECT 1814.770 101.220 1815.090 101.280 ;
        RECT 574.150 101.080 1815.090 101.220 ;
        RECT 574.150 101.020 574.470 101.080 ;
        RECT 1814.770 101.020 1815.090 101.080 ;
      LAYER via ;
        RECT 574.180 471.960 574.440 472.220 ;
        RECT 577.400 471.960 577.660 472.220 ;
        RECT 574.180 101.020 574.440 101.280 ;
        RECT 1814.800 101.020 1815.060 101.280 ;
      LAYER met2 ;
        RECT 577.650 500.000 577.930 504.000 ;
        RECT 577.690 498.850 577.830 500.000 ;
        RECT 577.460 498.710 577.830 498.850 ;
        RECT 577.460 472.250 577.600 498.710 ;
        RECT 574.180 471.930 574.440 472.250 ;
        RECT 577.400 471.930 577.660 472.250 ;
        RECT 574.240 101.310 574.380 471.930 ;
        RECT 574.180 100.990 574.440 101.310 ;
        RECT 1814.800 100.990 1815.060 101.310 ;
        RECT 1814.860 82.870 1815.000 100.990 ;
        RECT 1814.860 82.730 1817.760 82.870 ;
        RECT 1817.620 2.400 1817.760 82.730 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1829.030 16.900 1829.350 16.960 ;
        RECT 1835.010 16.900 1835.330 16.960 ;
        RECT 1829.030 16.760 1835.330 16.900 ;
        RECT 1829.030 16.700 1829.350 16.760 ;
        RECT 1835.010 16.700 1835.330 16.760 ;
      LAYER via ;
        RECT 1829.060 16.700 1829.320 16.960 ;
        RECT 1835.040 16.700 1835.300 16.960 ;
      LAYER met2 ;
        RECT 579.030 500.000 579.310 504.000 ;
        RECT 579.070 498.340 579.210 500.000 ;
        RECT 579.070 498.200 579.440 498.340 ;
        RECT 579.300 483.325 579.440 498.200 ;
        RECT 579.230 482.955 579.510 483.325 ;
        RECT 1829.050 65.435 1829.330 65.805 ;
        RECT 1829.120 16.990 1829.260 65.435 ;
        RECT 1829.060 16.670 1829.320 16.990 ;
        RECT 1835.040 16.670 1835.300 16.990 ;
        RECT 1835.100 2.400 1835.240 16.670 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
      LAYER via2 ;
        RECT 579.230 483.000 579.510 483.280 ;
        RECT 1829.050 65.480 1829.330 65.760 ;
      LAYER met3 ;
        RECT 579.205 483.300 579.535 483.305 ;
        RECT 578.950 483.290 579.535 483.300 ;
        RECT 578.750 482.990 579.535 483.290 ;
        RECT 578.950 482.980 579.535 482.990 ;
        RECT 579.205 482.975 579.535 482.980 ;
        RECT 578.950 65.770 579.330 65.780 ;
        RECT 1829.025 65.770 1829.355 65.785 ;
        RECT 578.950 65.470 1829.355 65.770 ;
        RECT 578.950 65.460 579.330 65.470 ;
        RECT 1829.025 65.455 1829.355 65.470 ;
      LAYER via3 ;
        RECT 578.980 482.980 579.300 483.300 ;
        RECT 578.980 65.460 579.300 65.780 ;
      LAYER met4 ;
        RECT 578.975 482.975 579.305 483.305 ;
        RECT 578.990 65.785 579.290 482.975 ;
        RECT 578.975 65.455 579.305 65.785 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.590 494.940 580.910 495.000 ;
        RECT 1849.270 494.940 1849.590 495.000 ;
        RECT 580.590 494.800 1849.590 494.940 ;
        RECT 580.590 494.740 580.910 494.800 ;
        RECT 1849.270 494.740 1849.590 494.800 ;
      LAYER via ;
        RECT 580.620 494.740 580.880 495.000 ;
        RECT 1849.300 494.740 1849.560 495.000 ;
      LAYER met2 ;
        RECT 580.410 500.000 580.690 504.000 ;
        RECT 580.450 499.360 580.590 500.000 ;
        RECT 580.450 499.220 580.820 499.360 ;
        RECT 580.680 495.030 580.820 499.220 ;
        RECT 580.620 494.710 580.880 495.030 ;
        RECT 1849.300 494.710 1849.560 495.030 ;
        RECT 1849.360 82.870 1849.500 494.710 ;
        RECT 1849.360 82.730 1850.880 82.870 ;
        RECT 1850.740 1.770 1850.880 82.730 ;
        RECT 1852.830 1.770 1853.390 2.400 ;
        RECT 1850.740 1.630 1853.390 1.770 ;
        RECT 1852.830 -4.800 1853.390 1.630 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.430 472.840 490.750 472.900 ;
        RECT 494.110 472.840 494.430 472.900 ;
        RECT 490.430 472.700 494.430 472.840 ;
        RECT 490.430 472.640 490.750 472.700 ;
        RECT 494.110 472.640 494.430 472.700 ;
        RECT 490.430 67.220 490.750 67.280 ;
        RECT 735.610 67.220 735.930 67.280 ;
        RECT 490.430 67.080 735.930 67.220 ;
        RECT 490.430 67.020 490.750 67.080 ;
        RECT 735.610 67.020 735.930 67.080 ;
      LAYER via ;
        RECT 490.460 472.640 490.720 472.900 ;
        RECT 494.140 472.640 494.400 472.900 ;
        RECT 490.460 67.020 490.720 67.280 ;
        RECT 735.640 67.020 735.900 67.280 ;
      LAYER met2 ;
        RECT 493.470 500.000 493.750 504.000 ;
        RECT 493.510 499.815 493.650 500.000 ;
        RECT 493.440 499.445 493.720 499.815 ;
        RECT 493.670 498.595 493.950 498.965 ;
        RECT 493.740 488.650 493.880 498.595 ;
        RECT 493.740 488.510 494.340 488.650 ;
        RECT 494.200 472.930 494.340 488.510 ;
        RECT 490.460 472.610 490.720 472.930 ;
        RECT 494.140 472.610 494.400 472.930 ;
        RECT 490.520 67.310 490.660 472.610 ;
        RECT 490.460 66.990 490.720 67.310 ;
        RECT 735.640 66.990 735.900 67.310 ;
        RECT 735.700 2.400 735.840 66.990 ;
        RECT 735.490 -4.800 736.050 2.400 ;
      LAYER via2 ;
        RECT 493.440 499.490 493.720 499.770 ;
        RECT 493.670 498.640 493.950 498.920 ;
      LAYER met3 ;
        RECT 493.415 499.465 493.745 499.795 ;
        RECT 493.430 498.945 493.730 499.465 ;
        RECT 493.430 498.630 493.975 498.945 ;
        RECT 493.645 498.615 493.975 498.630 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 581.510 109.040 581.830 109.100 ;
        RECT 1869.970 109.040 1870.290 109.100 ;
        RECT 581.510 108.900 1870.290 109.040 ;
        RECT 581.510 108.840 581.830 108.900 ;
        RECT 1869.970 108.840 1870.290 108.900 ;
      LAYER via ;
        RECT 581.540 108.840 581.800 109.100 ;
        RECT 1870.000 108.840 1870.260 109.100 ;
      LAYER met2 ;
        RECT 581.790 500.000 582.070 504.000 ;
        RECT 581.830 499.700 581.970 500.000 ;
        RECT 581.600 499.645 581.970 499.700 ;
        RECT 581.530 499.560 581.970 499.645 ;
        RECT 581.530 499.275 581.810 499.560 ;
        RECT 581.530 497.235 581.810 497.605 ;
        RECT 581.600 109.130 581.740 497.235 ;
        RECT 581.540 108.810 581.800 109.130 ;
        RECT 1870.000 108.810 1870.260 109.130 ;
        RECT 1870.060 5.850 1870.200 108.810 ;
        RECT 1870.060 5.710 1870.660 5.850 ;
        RECT 1870.520 2.400 1870.660 5.710 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
      LAYER via2 ;
        RECT 581.530 499.320 581.810 499.600 ;
        RECT 581.530 497.280 581.810 497.560 ;
      LAYER met3 ;
        RECT 581.505 499.610 581.835 499.625 ;
        RECT 581.505 499.295 582.050 499.610 ;
        RECT 581.750 497.585 582.050 499.295 ;
        RECT 581.505 497.270 582.050 497.585 ;
        RECT 581.505 497.255 581.835 497.270 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.130 491.540 580.450 491.600 ;
        RECT 582.890 491.540 583.210 491.600 ;
        RECT 580.130 491.400 583.210 491.540 ;
        RECT 580.130 491.340 580.450 491.400 ;
        RECT 582.890 491.340 583.210 491.400 ;
        RECT 579.670 45.460 579.990 45.520 ;
        RECT 1888.370 45.460 1888.690 45.520 ;
        RECT 579.670 45.320 1888.690 45.460 ;
        RECT 579.670 45.260 579.990 45.320 ;
        RECT 1888.370 45.260 1888.690 45.320 ;
      LAYER via ;
        RECT 580.160 491.340 580.420 491.600 ;
        RECT 582.920 491.340 583.180 491.600 ;
        RECT 579.700 45.260 579.960 45.520 ;
        RECT 1888.400 45.260 1888.660 45.520 ;
      LAYER met2 ;
        RECT 583.170 500.000 583.450 504.000 ;
        RECT 583.210 498.680 583.350 500.000 ;
        RECT 582.980 498.540 583.350 498.680 ;
        RECT 582.980 491.630 583.120 498.540 ;
        RECT 580.160 491.310 580.420 491.630 ;
        RECT 582.920 491.310 583.180 491.630 ;
        RECT 580.220 473.010 580.360 491.310 ;
        RECT 579.760 472.870 580.360 473.010 ;
        RECT 579.760 45.550 579.900 472.870 ;
        RECT 579.700 45.230 579.960 45.550 ;
        RECT 1888.400 45.230 1888.660 45.550 ;
        RECT 1888.460 2.400 1888.600 45.230 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 584.500 499.500 584.820 499.760 ;
        RECT 584.590 499.080 584.730 499.500 ;
        RECT 584.590 498.880 585.050 499.080 ;
        RECT 584.730 498.820 585.050 498.880 ;
      LAYER via ;
        RECT 584.530 499.500 584.790 499.760 ;
        RECT 584.760 498.820 585.020 499.080 ;
      LAYER met2 ;
        RECT 584.550 500.000 584.830 504.000 ;
        RECT 584.590 499.790 584.730 500.000 ;
        RECT 584.530 499.470 584.790 499.790 ;
        RECT 584.760 498.965 585.020 499.110 ;
        RECT 584.750 498.595 585.030 498.965 ;
        RECT 1905.870 64.755 1906.150 65.125 ;
        RECT 1905.940 2.400 1906.080 64.755 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
      LAYER via2 ;
        RECT 584.750 498.640 585.030 498.920 ;
        RECT 1905.870 64.800 1906.150 65.080 ;
      LAYER met3 ;
        RECT 584.725 498.930 585.055 498.945 ;
        RECT 585.390 498.930 585.770 498.940 ;
        RECT 584.725 498.630 585.770 498.930 ;
        RECT 584.725 498.615 585.055 498.630 ;
        RECT 585.390 498.620 585.770 498.630 ;
        RECT 585.390 65.090 585.770 65.100 ;
        RECT 1905.845 65.090 1906.175 65.105 ;
        RECT 585.390 64.790 1906.175 65.090 ;
        RECT 585.390 64.780 585.770 64.790 ;
        RECT 1905.845 64.775 1906.175 64.790 ;
      LAYER via3 ;
        RECT 585.420 498.620 585.740 498.940 ;
        RECT 585.420 64.780 585.740 65.100 ;
      LAYER met4 ;
        RECT 585.415 498.615 585.745 498.945 ;
        RECT 585.430 65.105 585.730 498.615 ;
        RECT 585.415 64.775 585.745 65.105 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.930 500.000 586.210 504.000 ;
        RECT 585.970 498.680 586.110 500.000 ;
        RECT 585.970 498.540 586.340 498.680 ;
        RECT 586.200 489.445 586.340 498.540 ;
        RECT 586.130 489.075 586.410 489.445 ;
        RECT 1921.510 72.915 1921.790 73.285 ;
        RECT 1921.580 1.770 1921.720 72.915 ;
        RECT 1923.670 1.770 1924.230 2.400 ;
        RECT 1921.580 1.630 1924.230 1.770 ;
        RECT 1923.670 -4.800 1924.230 1.630 ;
      LAYER via2 ;
        RECT 586.130 489.120 586.410 489.400 ;
        RECT 1921.510 72.960 1921.790 73.240 ;
      LAYER met3 ;
        RECT 584.470 489.410 584.850 489.420 ;
        RECT 586.105 489.410 586.435 489.425 ;
        RECT 584.470 489.110 586.435 489.410 ;
        RECT 584.470 489.100 584.850 489.110 ;
        RECT 586.105 489.095 586.435 489.110 ;
        RECT 584.470 73.250 584.850 73.260 ;
        RECT 1921.485 73.250 1921.815 73.265 ;
        RECT 584.470 72.950 1921.815 73.250 ;
        RECT 584.470 72.940 584.850 72.950 ;
        RECT 1921.485 72.935 1921.815 72.950 ;
      LAYER via3 ;
        RECT 584.500 489.100 584.820 489.420 ;
        RECT 584.500 72.940 584.820 73.260 ;
      LAYER met4 ;
        RECT 584.495 489.095 584.825 489.425 ;
        RECT 584.510 73.265 584.810 489.095 ;
        RECT 584.495 72.935 584.825 73.265 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.730 494.600 608.050 494.660 ;
        RECT 1938.970 494.600 1939.290 494.660 ;
        RECT 607.730 494.460 1939.290 494.600 ;
        RECT 607.730 494.400 608.050 494.460 ;
        RECT 1938.970 494.400 1939.290 494.460 ;
      LAYER via ;
        RECT 607.760 494.400 608.020 494.660 ;
        RECT 1939.000 494.400 1939.260 494.660 ;
      LAYER met2 ;
        RECT 587.310 500.000 587.590 504.000 ;
        RECT 587.350 499.020 587.490 500.000 ;
        RECT 587.120 498.880 587.490 499.020 ;
        RECT 587.120 495.565 587.260 498.880 ;
        RECT 587.050 495.195 587.330 495.565 ;
        RECT 607.750 495.195 608.030 495.565 ;
        RECT 607.820 494.690 607.960 495.195 ;
        RECT 607.760 494.370 608.020 494.690 ;
        RECT 1939.000 494.370 1939.260 494.690 ;
        RECT 1939.060 1.770 1939.200 494.370 ;
        RECT 1941.150 1.770 1941.710 2.400 ;
        RECT 1939.060 1.630 1941.710 1.770 ;
        RECT 1941.150 -4.800 1941.710 1.630 ;
      LAYER via2 ;
        RECT 587.050 495.240 587.330 495.520 ;
        RECT 607.750 495.240 608.030 495.520 ;
      LAYER met3 ;
        RECT 587.025 495.530 587.355 495.545 ;
        RECT 607.725 495.530 608.055 495.545 ;
        RECT 587.025 495.230 608.055 495.530 ;
        RECT 587.025 495.215 587.355 495.230 ;
        RECT 607.725 495.215 608.055 495.230 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 588.410 108.360 588.730 108.420 ;
        RECT 1952.770 108.360 1953.090 108.420 ;
        RECT 588.410 108.220 1953.090 108.360 ;
        RECT 588.410 108.160 588.730 108.220 ;
        RECT 1952.770 108.160 1953.090 108.220 ;
        RECT 1952.770 16.900 1953.090 16.960 ;
        RECT 1959.210 16.900 1959.530 16.960 ;
        RECT 1952.770 16.760 1959.530 16.900 ;
        RECT 1952.770 16.700 1953.090 16.760 ;
        RECT 1959.210 16.700 1959.530 16.760 ;
      LAYER via ;
        RECT 588.440 108.160 588.700 108.420 ;
        RECT 1952.800 108.160 1953.060 108.420 ;
        RECT 1952.800 16.700 1953.060 16.960 ;
        RECT 1959.240 16.700 1959.500 16.960 ;
      LAYER met2 ;
        RECT 588.690 500.000 588.970 504.000 ;
        RECT 588.730 498.850 588.870 500.000 ;
        RECT 588.500 498.710 588.870 498.850 ;
        RECT 588.500 108.450 588.640 498.710 ;
        RECT 588.440 108.130 588.700 108.450 ;
        RECT 1952.800 108.130 1953.060 108.450 ;
        RECT 1952.860 16.990 1953.000 108.130 ;
        RECT 1952.800 16.670 1953.060 16.990 ;
        RECT 1959.240 16.670 1959.500 16.990 ;
        RECT 1959.300 2.400 1959.440 16.670 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 590.020 499.500 590.340 499.760 ;
        RECT 590.110 498.060 590.250 499.500 ;
        RECT 589.790 497.860 590.250 498.060 ;
        RECT 589.790 497.800 590.110 497.860 ;
        RECT 587.950 491.540 588.270 491.600 ;
        RECT 589.790 491.540 590.110 491.600 ;
        RECT 587.950 491.400 590.110 491.540 ;
        RECT 587.950 491.340 588.270 491.400 ;
        RECT 589.790 491.340 590.110 491.400 ;
        RECT 587.950 108.020 588.270 108.080 ;
        RECT 1973.470 108.020 1973.790 108.080 ;
        RECT 587.950 107.880 1973.790 108.020 ;
        RECT 587.950 107.820 588.270 107.880 ;
        RECT 1973.470 107.820 1973.790 107.880 ;
      LAYER via ;
        RECT 590.050 499.500 590.310 499.760 ;
        RECT 589.820 497.800 590.080 498.060 ;
        RECT 587.980 491.340 588.240 491.600 ;
        RECT 589.820 491.340 590.080 491.600 ;
        RECT 587.980 107.820 588.240 108.080 ;
        RECT 1973.500 107.820 1973.760 108.080 ;
      LAYER met2 ;
        RECT 590.070 500.000 590.350 504.000 ;
        RECT 590.110 499.790 590.250 500.000 ;
        RECT 590.050 499.470 590.310 499.790 ;
        RECT 589.820 497.770 590.080 498.090 ;
        RECT 589.880 491.630 590.020 497.770 ;
        RECT 587.980 491.310 588.240 491.630 ;
        RECT 589.820 491.310 590.080 491.630 ;
        RECT 588.040 108.110 588.180 491.310 ;
        RECT 587.980 107.790 588.240 108.110 ;
        RECT 1973.500 107.790 1973.760 108.110 ;
        RECT 1973.560 82.870 1973.700 107.790 ;
        RECT 1973.560 82.730 1976.920 82.870 ;
        RECT 1976.780 2.400 1976.920 82.730 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.450 500.000 591.730 504.000 ;
        RECT 591.490 499.645 591.630 500.000 ;
        RECT 591.420 499.275 591.700 499.645 ;
        RECT 1994.650 72.235 1994.930 72.605 ;
        RECT 1994.720 2.400 1994.860 72.235 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
      LAYER via2 ;
        RECT 591.420 499.320 591.700 499.600 ;
        RECT 1994.650 72.280 1994.930 72.560 ;
      LAYER met3 ;
        RECT 591.395 499.610 591.725 499.625 ;
        RECT 592.750 499.610 593.130 499.620 ;
        RECT 591.395 499.310 593.130 499.610 ;
        RECT 591.395 499.295 591.725 499.310 ;
        RECT 592.750 499.300 593.130 499.310 ;
        RECT 592.750 72.570 593.130 72.580 ;
        RECT 1994.625 72.570 1994.955 72.585 ;
        RECT 592.750 72.270 1994.955 72.570 ;
        RECT 592.750 72.260 593.130 72.270 ;
        RECT 1994.625 72.255 1994.955 72.270 ;
      LAYER via3 ;
        RECT 592.780 499.300 593.100 499.620 ;
        RECT 592.780 72.260 593.100 72.580 ;
      LAYER met4 ;
        RECT 592.775 499.295 593.105 499.625 ;
        RECT 592.790 72.585 593.090 499.295 ;
        RECT 592.775 72.255 593.105 72.585 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 592.780 499.500 593.100 499.760 ;
        RECT 592.870 498.400 593.010 499.500 ;
        RECT 592.870 498.200 593.330 498.400 ;
        RECT 593.010 498.140 593.330 498.200 ;
      LAYER via ;
        RECT 592.810 499.500 593.070 499.760 ;
        RECT 593.040 498.140 593.300 498.400 ;
      LAYER met2 ;
        RECT 592.830 500.000 593.110 504.000 ;
        RECT 592.870 499.790 593.010 500.000 ;
        RECT 592.810 499.470 593.070 499.790 ;
        RECT 593.040 498.110 593.300 498.430 ;
        RECT 593.100 494.885 593.240 498.110 ;
        RECT 593.030 494.515 593.310 494.885 ;
        RECT 2012.590 79.715 2012.870 80.085 ;
        RECT 2012.660 2.400 2012.800 79.715 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
      LAYER via2 ;
        RECT 593.030 494.560 593.310 494.840 ;
        RECT 2012.590 79.760 2012.870 80.040 ;
      LAYER met3 ;
        RECT 591.830 494.850 592.210 494.860 ;
        RECT 593.005 494.850 593.335 494.865 ;
        RECT 591.830 494.550 593.335 494.850 ;
        RECT 591.830 494.540 592.210 494.550 ;
        RECT 593.005 494.535 593.335 494.550 ;
        RECT 591.830 80.050 592.210 80.060 ;
        RECT 2012.565 80.050 2012.895 80.065 ;
        RECT 591.830 79.750 2012.895 80.050 ;
        RECT 591.830 79.740 592.210 79.750 ;
        RECT 2012.565 79.735 2012.895 79.750 ;
      LAYER via3 ;
        RECT 591.860 494.540 592.180 494.860 ;
        RECT 591.860 79.740 592.180 80.060 ;
      LAYER met4 ;
        RECT 591.855 494.535 592.185 494.865 ;
        RECT 591.870 80.065 592.170 494.535 ;
        RECT 591.855 79.735 592.185 80.065 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.390 493.920 594.710 493.980 ;
        RECT 2028.670 493.920 2028.990 493.980 ;
        RECT 594.390 493.780 2028.990 493.920 ;
        RECT 594.390 493.720 594.710 493.780 ;
        RECT 2028.670 493.720 2028.990 493.780 ;
      LAYER via ;
        RECT 594.420 493.720 594.680 493.980 ;
        RECT 2028.700 493.720 2028.960 493.980 ;
      LAYER met2 ;
        RECT 594.210 500.000 594.490 504.000 ;
        RECT 594.250 498.340 594.390 500.000 ;
        RECT 594.250 498.200 594.620 498.340 ;
        RECT 594.480 494.010 594.620 498.200 ;
        RECT 594.420 493.690 594.680 494.010 ;
        RECT 2028.700 493.690 2028.960 494.010 ;
        RECT 2028.760 82.870 2028.900 493.690 ;
        RECT 2028.760 82.730 2030.280 82.870 ;
        RECT 2030.140 2.400 2030.280 82.730 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 494.800 499.700 495.120 499.760 ;
        RECT 494.800 499.500 495.260 499.700 ;
        RECT 495.120 498.400 495.260 499.500 ;
        RECT 495.030 498.140 495.350 498.400 ;
      LAYER via ;
        RECT 494.830 499.500 495.090 499.760 ;
        RECT 495.060 498.140 495.320 498.400 ;
      LAYER met2 ;
        RECT 494.850 500.000 495.130 504.000 ;
        RECT 494.890 499.790 495.030 500.000 ;
        RECT 494.830 499.470 495.090 499.790 ;
        RECT 495.060 498.285 495.320 498.430 ;
        RECT 495.050 497.915 495.330 498.285 ;
        RECT 753.110 78.355 753.390 78.725 ;
        RECT 753.180 2.400 753.320 78.355 ;
        RECT 752.970 -4.800 753.530 2.400 ;
      LAYER via2 ;
        RECT 495.050 497.960 495.330 498.240 ;
        RECT 753.110 78.400 753.390 78.680 ;
      LAYER met3 ;
        RECT 495.025 498.250 495.355 498.265 ;
        RECT 496.150 498.250 496.530 498.260 ;
        RECT 495.025 497.950 496.530 498.250 ;
        RECT 495.025 497.935 495.355 497.950 ;
        RECT 496.150 497.940 496.530 497.950 ;
        RECT 496.150 78.690 496.530 78.700 ;
        RECT 753.085 78.690 753.415 78.705 ;
        RECT 496.150 78.390 753.415 78.690 ;
        RECT 496.150 78.380 496.530 78.390 ;
        RECT 753.085 78.375 753.415 78.390 ;
      LAYER via3 ;
        RECT 496.180 497.940 496.500 498.260 ;
        RECT 496.180 78.380 496.500 78.700 ;
      LAYER met4 ;
        RECT 496.175 497.935 496.505 498.265 ;
        RECT 496.190 78.705 496.490 497.935 ;
        RECT 496.175 78.375 496.505 78.705 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 595.310 474.000 595.630 474.260 ;
        RECT 595.400 473.240 595.540 474.000 ;
        RECT 595.310 472.980 595.630 473.240 ;
        RECT 595.310 115.840 595.630 115.900 ;
        RECT 2042.470 115.840 2042.790 115.900 ;
        RECT 595.310 115.700 2042.790 115.840 ;
        RECT 595.310 115.640 595.630 115.700 ;
        RECT 2042.470 115.640 2042.790 115.700 ;
      LAYER via ;
        RECT 595.340 474.000 595.600 474.260 ;
        RECT 595.340 472.980 595.600 473.240 ;
        RECT 595.340 115.640 595.600 115.900 ;
        RECT 2042.500 115.640 2042.760 115.900 ;
      LAYER met2 ;
        RECT 595.590 500.000 595.870 504.000 ;
        RECT 595.630 499.815 595.770 500.000 ;
        RECT 595.560 499.445 595.840 499.815 ;
        RECT 595.330 494.515 595.610 494.885 ;
        RECT 595.400 474.290 595.540 494.515 ;
        RECT 595.340 473.970 595.600 474.290 ;
        RECT 595.340 472.950 595.600 473.270 ;
        RECT 595.400 115.930 595.540 472.950 ;
        RECT 595.340 115.610 595.600 115.930 ;
        RECT 2042.500 115.610 2042.760 115.930 ;
        RECT 2042.560 82.870 2042.700 115.610 ;
        RECT 2042.560 82.730 2045.920 82.870 ;
        RECT 2045.780 1.770 2045.920 82.730 ;
        RECT 2047.870 1.770 2048.430 2.400 ;
        RECT 2045.780 1.630 2048.430 1.770 ;
        RECT 2047.870 -4.800 2048.430 1.630 ;
      LAYER via2 ;
        RECT 595.560 499.490 595.840 499.770 ;
        RECT 595.330 494.560 595.610 494.840 ;
      LAYER met3 ;
        RECT 595.535 499.620 595.865 499.795 ;
        RECT 595.510 499.610 595.890 499.620 ;
        RECT 595.510 499.310 596.150 499.610 ;
        RECT 595.510 499.300 595.890 499.310 ;
        RECT 595.305 494.860 595.635 494.865 ;
        RECT 595.305 494.850 595.890 494.860 ;
        RECT 595.080 494.550 595.890 494.850 ;
        RECT 595.305 494.540 595.890 494.550 ;
        RECT 595.305 494.535 595.635 494.540 ;
      LAYER via3 ;
        RECT 595.540 499.300 595.860 499.620 ;
        RECT 595.540 494.540 595.860 494.860 ;
      LAYER met4 ;
        RECT 595.535 499.295 595.865 499.625 ;
        RECT 595.550 494.865 595.850 499.295 ;
        RECT 595.535 494.535 595.865 494.865 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 596.920 499.700 597.240 499.760 ;
        RECT 596.550 499.560 597.240 499.700 ;
        RECT 596.550 498.740 596.690 499.560 ;
        RECT 596.920 499.500 597.240 499.560 ;
        RECT 596.230 498.540 596.690 498.740 ;
        RECT 596.230 498.480 596.550 498.540 ;
        RECT 594.850 115.500 595.170 115.560 ;
        RECT 2063.170 115.500 2063.490 115.560 ;
        RECT 594.850 115.360 2063.490 115.500 ;
        RECT 594.850 115.300 595.170 115.360 ;
        RECT 2063.170 115.300 2063.490 115.360 ;
      LAYER via ;
        RECT 596.950 499.500 597.210 499.760 ;
        RECT 596.260 498.480 596.520 498.740 ;
        RECT 594.880 115.300 595.140 115.560 ;
        RECT 2063.200 115.300 2063.460 115.560 ;
      LAYER met2 ;
        RECT 596.970 500.000 597.250 504.000 ;
        RECT 597.010 499.790 597.150 500.000 ;
        RECT 596.950 499.470 597.210 499.790 ;
        RECT 596.260 498.450 596.520 498.770 ;
        RECT 596.320 473.690 596.460 498.450 ;
        RECT 594.940 473.550 596.460 473.690 ;
        RECT 594.940 115.590 595.080 473.550 ;
        RECT 594.880 115.270 595.140 115.590 ;
        RECT 2063.200 115.270 2063.460 115.590 ;
        RECT 2063.260 1.770 2063.400 115.270 ;
        RECT 2065.350 1.770 2065.910 2.400 ;
        RECT 2063.260 1.630 2065.910 1.770 ;
        RECT 2065.350 -4.800 2065.910 1.630 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 598.300 499.500 598.620 499.760 ;
        RECT 598.390 498.000 598.530 499.500 ;
        RECT 598.990 498.000 599.310 498.060 ;
        RECT 598.390 497.860 599.310 498.000 ;
        RECT 598.990 497.800 599.310 497.860 ;
        RECT 593.930 466.720 594.250 466.780 ;
        RECT 598.070 466.720 598.390 466.780 ;
        RECT 593.930 466.580 598.390 466.720 ;
        RECT 593.930 466.520 594.250 466.580 ;
        RECT 598.070 466.520 598.390 466.580 ;
        RECT 593.930 86.600 594.250 86.660 ;
        RECT 2077.430 86.600 2077.750 86.660 ;
        RECT 593.930 86.460 2077.750 86.600 ;
        RECT 593.930 86.400 594.250 86.460 ;
        RECT 2077.430 86.400 2077.750 86.460 ;
        RECT 2077.430 16.900 2077.750 16.960 ;
        RECT 2083.410 16.900 2083.730 16.960 ;
        RECT 2077.430 16.760 2083.730 16.900 ;
        RECT 2077.430 16.700 2077.750 16.760 ;
        RECT 2083.410 16.700 2083.730 16.760 ;
      LAYER via ;
        RECT 598.330 499.500 598.590 499.760 ;
        RECT 599.020 497.800 599.280 498.060 ;
        RECT 593.960 466.520 594.220 466.780 ;
        RECT 598.100 466.520 598.360 466.780 ;
        RECT 593.960 86.400 594.220 86.660 ;
        RECT 2077.460 86.400 2077.720 86.660 ;
        RECT 2077.460 16.700 2077.720 16.960 ;
        RECT 2083.440 16.700 2083.700 16.960 ;
      LAYER met2 ;
        RECT 598.350 500.000 598.630 504.000 ;
        RECT 598.390 499.790 598.530 500.000 ;
        RECT 598.330 499.470 598.590 499.790 ;
        RECT 599.020 497.770 599.280 498.090 ;
        RECT 599.080 489.970 599.220 497.770 ;
        RECT 598.620 489.830 599.220 489.970 ;
        RECT 598.620 483.070 598.760 489.830 ;
        RECT 598.160 482.930 598.760 483.070 ;
        RECT 598.160 466.810 598.300 482.930 ;
        RECT 593.960 466.490 594.220 466.810 ;
        RECT 598.100 466.490 598.360 466.810 ;
        RECT 594.020 86.690 594.160 466.490 ;
        RECT 593.960 86.370 594.220 86.690 ;
        RECT 2077.460 86.370 2077.720 86.690 ;
        RECT 2077.520 16.990 2077.660 86.370 ;
        RECT 2077.460 16.670 2077.720 16.990 ;
        RECT 2083.440 16.670 2083.700 16.990 ;
        RECT 2083.500 2.400 2083.640 16.670 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.730 500.000 600.010 504.000 ;
        RECT 599.770 499.645 599.910 500.000 ;
        RECT 599.700 499.275 599.980 499.645 ;
        RECT 2097.690 85.835 2097.970 86.205 ;
        RECT 2097.760 82.870 2097.900 85.835 ;
        RECT 2097.760 82.730 2101.120 82.870 ;
        RECT 2100.980 2.400 2101.120 82.730 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
      LAYER via2 ;
        RECT 599.700 499.320 599.980 499.600 ;
        RECT 2097.690 85.880 2097.970 86.160 ;
      LAYER met3 ;
        RECT 599.190 500.290 599.570 500.300 ;
        RECT 599.000 499.980 599.570 500.290 ;
        RECT 599.000 499.610 599.300 499.980 ;
        RECT 599.675 499.610 600.005 499.625 ;
        RECT 599.000 499.310 600.005 499.610 ;
        RECT 599.675 499.295 600.005 499.310 ;
        RECT 599.190 86.170 599.570 86.180 ;
        RECT 2097.665 86.170 2097.995 86.185 ;
        RECT 599.190 85.870 2097.995 86.170 ;
        RECT 599.190 85.860 599.570 85.870 ;
        RECT 2097.665 85.855 2097.995 85.870 ;
      LAYER via3 ;
        RECT 599.220 499.980 599.540 500.300 ;
        RECT 599.220 85.860 599.540 86.180 ;
      LAYER met4 ;
        RECT 599.215 499.975 599.545 500.305 ;
        RECT 599.230 86.185 599.530 499.975 ;
        RECT 599.215 85.855 599.545 86.185 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 601.150 499.900 604.050 500.040 ;
        RECT 601.150 499.760 601.290 499.900 ;
        RECT 601.060 499.500 601.380 499.760 ;
        RECT 603.910 497.660 604.050 499.900 ;
        RECT 605.890 497.660 606.210 497.720 ;
        RECT 603.910 497.520 606.210 497.660 ;
        RECT 605.890 497.460 606.210 497.520 ;
        RECT 605.890 493.580 606.210 493.640 ;
        RECT 2118.370 493.580 2118.690 493.640 ;
        RECT 605.890 493.440 2118.690 493.580 ;
        RECT 605.890 493.380 606.210 493.440 ;
        RECT 2118.370 493.380 2118.690 493.440 ;
      LAYER via ;
        RECT 601.090 499.500 601.350 499.760 ;
        RECT 605.920 497.460 606.180 497.720 ;
        RECT 605.920 493.380 606.180 493.640 ;
        RECT 2118.400 493.380 2118.660 493.640 ;
      LAYER met2 ;
        RECT 601.110 500.000 601.390 504.000 ;
        RECT 601.150 499.790 601.290 500.000 ;
        RECT 601.090 499.470 601.350 499.790 ;
        RECT 605.920 497.430 606.180 497.750 ;
        RECT 605.980 493.670 606.120 497.430 ;
        RECT 605.920 493.350 606.180 493.670 ;
        RECT 2118.400 493.350 2118.660 493.670 ;
        RECT 2118.460 16.050 2118.600 493.350 ;
        RECT 2118.460 15.910 2119.060 16.050 ;
        RECT 2118.920 2.400 2119.060 15.910 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 601.290 496.980 601.610 497.040 ;
        RECT 602.210 496.980 602.530 497.040 ;
        RECT 601.290 496.840 602.530 496.980 ;
        RECT 601.290 496.780 601.610 496.840 ;
        RECT 602.210 496.780 602.530 496.840 ;
        RECT 601.290 115.160 601.610 115.220 ;
        RECT 2132.170 115.160 2132.490 115.220 ;
        RECT 601.290 115.020 2132.490 115.160 ;
        RECT 601.290 114.960 601.610 115.020 ;
        RECT 2132.170 114.960 2132.490 115.020 ;
      LAYER via ;
        RECT 601.320 496.780 601.580 497.040 ;
        RECT 602.240 496.780 602.500 497.040 ;
        RECT 601.320 114.960 601.580 115.220 ;
        RECT 2132.200 114.960 2132.460 115.220 ;
      LAYER met2 ;
        RECT 602.490 500.000 602.770 504.000 ;
        RECT 602.530 498.850 602.670 500.000 ;
        RECT 602.300 498.710 602.670 498.850 ;
        RECT 602.300 497.070 602.440 498.710 ;
        RECT 601.320 496.750 601.580 497.070 ;
        RECT 602.240 496.750 602.500 497.070 ;
        RECT 601.380 115.250 601.520 496.750 ;
        RECT 601.320 114.930 601.580 115.250 ;
        RECT 2132.200 114.930 2132.460 115.250 ;
        RECT 2132.260 82.870 2132.400 114.930 ;
        RECT 2132.260 82.730 2134.240 82.870 ;
        RECT 2134.100 1.770 2134.240 82.730 ;
        RECT 2136.190 1.770 2136.750 2.400 ;
        RECT 2134.100 1.630 2136.750 1.770 ;
        RECT 2136.190 -4.800 2136.750 1.630 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.830 462.980 601.150 463.040 ;
        RECT 603.590 462.980 603.910 463.040 ;
        RECT 600.830 462.840 603.910 462.980 ;
        RECT 600.830 462.780 601.150 462.840 ;
        RECT 603.590 462.780 603.910 462.840 ;
        RECT 600.830 114.480 601.150 114.540 ;
        RECT 2152.870 114.480 2153.190 114.540 ;
        RECT 600.830 114.340 2153.190 114.480 ;
        RECT 600.830 114.280 601.150 114.340 ;
        RECT 2152.870 114.280 2153.190 114.340 ;
      LAYER via ;
        RECT 600.860 462.780 601.120 463.040 ;
        RECT 603.620 462.780 603.880 463.040 ;
        RECT 600.860 114.280 601.120 114.540 ;
        RECT 2152.900 114.280 2153.160 114.540 ;
      LAYER met2 ;
        RECT 603.870 500.000 604.150 504.000 ;
        RECT 603.910 499.815 604.050 500.000 ;
        RECT 603.840 499.445 604.120 499.815 ;
        RECT 603.610 498.595 603.890 498.965 ;
        RECT 603.680 463.070 603.820 498.595 ;
        RECT 600.860 462.750 601.120 463.070 ;
        RECT 603.620 462.750 603.880 463.070 ;
        RECT 600.920 114.570 601.060 462.750 ;
        RECT 600.860 114.250 601.120 114.570 ;
        RECT 2152.900 114.250 2153.160 114.570 ;
        RECT 2152.960 82.870 2153.100 114.250 ;
        RECT 2152.960 82.730 2154.480 82.870 ;
        RECT 2154.340 2.400 2154.480 82.730 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
      LAYER via2 ;
        RECT 603.840 499.490 604.120 499.770 ;
        RECT 603.610 498.640 603.890 498.920 ;
      LAYER met3 ;
        RECT 603.815 499.465 604.145 499.795 ;
        RECT 603.830 498.945 604.130 499.465 ;
        RECT 603.585 498.630 604.130 498.945 ;
        RECT 603.585 498.615 603.915 498.630 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.250 500.000 605.530 504.000 ;
        RECT 605.290 498.965 605.430 500.000 ;
        RECT 605.220 498.595 605.500 498.965 ;
        RECT 2166.690 93.995 2166.970 94.365 ;
        RECT 2166.760 82.870 2166.900 93.995 ;
        RECT 2166.760 82.730 2170.120 82.870 ;
        RECT 2169.980 1.770 2170.120 82.730 ;
        RECT 2172.070 1.770 2172.630 2.400 ;
        RECT 2169.980 1.630 2172.630 1.770 ;
        RECT 2172.070 -4.800 2172.630 1.630 ;
      LAYER via2 ;
        RECT 605.220 498.640 605.500 498.920 ;
        RECT 2166.690 94.040 2166.970 94.320 ;
      LAYER met3 ;
        RECT 605.195 498.930 605.525 498.945 ;
        RECT 605.195 498.615 605.740 498.930 ;
        RECT 605.440 498.260 605.740 498.615 ;
        RECT 605.440 497.950 606.010 498.260 ;
        RECT 605.630 497.940 606.010 497.950 ;
        RECT 605.630 94.330 606.010 94.340 ;
        RECT 2166.665 94.330 2166.995 94.345 ;
        RECT 605.630 94.030 2166.995 94.330 ;
        RECT 605.630 94.020 606.010 94.030 ;
        RECT 2166.665 94.015 2166.995 94.030 ;
      LAYER via3 ;
        RECT 605.660 497.940 605.980 498.260 ;
        RECT 605.660 94.020 605.980 94.340 ;
      LAYER met4 ;
        RECT 605.655 497.935 605.985 498.265 ;
        RECT 605.670 94.345 605.970 497.935 ;
        RECT 605.655 94.015 605.985 94.345 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.630 500.000 606.910 504.000 ;
        RECT 606.670 499.815 606.810 500.000 ;
        RECT 606.600 499.445 606.880 499.815 ;
        RECT 2187.390 93.315 2187.670 93.685 ;
        RECT 2187.460 1.770 2187.600 93.315 ;
        RECT 2189.550 1.770 2190.110 2.400 ;
        RECT 2187.460 1.630 2190.110 1.770 ;
        RECT 2189.550 -4.800 2190.110 1.630 ;
      LAYER via2 ;
        RECT 606.600 499.490 606.880 499.770 ;
        RECT 2187.390 93.360 2187.670 93.640 ;
      LAYER met3 ;
        RECT 606.575 499.620 606.905 499.795 ;
        RECT 606.550 499.610 606.930 499.620 ;
        RECT 606.550 499.310 607.190 499.610 ;
        RECT 606.550 499.300 606.930 499.310 ;
        RECT 606.550 93.650 606.930 93.660 ;
        RECT 2187.365 93.650 2187.695 93.665 ;
        RECT 606.550 93.350 2187.695 93.650 ;
        RECT 606.550 93.340 606.930 93.350 ;
        RECT 2187.365 93.335 2187.695 93.350 ;
      LAYER via3 ;
        RECT 606.580 499.300 606.900 499.620 ;
        RECT 606.580 93.340 606.900 93.660 ;
      LAYER met4 ;
        RECT 606.575 499.295 606.905 499.625 ;
        RECT 606.590 93.665 606.890 499.295 ;
        RECT 606.575 93.335 606.905 93.665 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 665.690 501.740 666.010 501.800 ;
        RECT 607.130 501.600 666.010 501.740 ;
        RECT 607.130 499.360 607.270 501.600 ;
        RECT 665.690 501.540 666.010 501.600 ;
        RECT 607.960 499.360 608.280 499.420 ;
        RECT 607.130 499.220 608.280 499.360 ;
        RECT 607.960 499.160 608.280 499.220 ;
        RECT 665.690 497.660 666.010 497.720 ;
        RECT 2201.170 497.660 2201.490 497.720 ;
        RECT 665.690 497.520 2201.490 497.660 ;
        RECT 665.690 497.460 666.010 497.520 ;
        RECT 2201.170 497.460 2201.490 497.520 ;
        RECT 2201.170 16.900 2201.490 16.960 ;
        RECT 2207.610 16.900 2207.930 16.960 ;
        RECT 2201.170 16.760 2207.930 16.900 ;
        RECT 2201.170 16.700 2201.490 16.760 ;
        RECT 2207.610 16.700 2207.930 16.760 ;
      LAYER via ;
        RECT 665.720 501.540 665.980 501.800 ;
        RECT 607.990 499.160 608.250 499.420 ;
        RECT 665.720 497.460 665.980 497.720 ;
        RECT 2201.200 497.460 2201.460 497.720 ;
        RECT 2201.200 16.700 2201.460 16.960 ;
        RECT 2207.640 16.700 2207.900 16.960 ;
      LAYER met2 ;
        RECT 608.010 500.000 608.290 504.000 ;
        RECT 665.720 501.510 665.980 501.830 ;
        RECT 608.050 499.450 608.190 500.000 ;
        RECT 607.990 499.130 608.250 499.450 ;
        RECT 665.780 497.750 665.920 501.510 ;
        RECT 665.720 497.430 665.980 497.750 ;
        RECT 2201.200 497.430 2201.460 497.750 ;
        RECT 2201.260 16.990 2201.400 497.430 ;
        RECT 2201.200 16.670 2201.460 16.990 ;
        RECT 2207.640 16.670 2207.900 16.990 ;
        RECT 2207.700 2.400 2207.840 16.670 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.230 500.000 496.510 504.000 ;
        RECT 496.270 498.340 496.410 500.000 ;
        RECT 496.270 498.200 496.640 498.340 ;
        RECT 496.500 485.365 496.640 498.200 ;
        RECT 496.430 484.995 496.710 485.365 ;
        RECT 765.990 121.875 766.270 122.245 ;
        RECT 766.060 82.870 766.200 121.875 ;
        RECT 766.060 82.730 768.960 82.870 ;
        RECT 768.820 1.770 768.960 82.730 ;
        RECT 770.910 1.770 771.470 2.400 ;
        RECT 768.820 1.630 771.470 1.770 ;
        RECT 770.910 -4.800 771.470 1.630 ;
      LAYER via2 ;
        RECT 496.430 485.040 496.710 485.320 ;
        RECT 765.990 121.920 766.270 122.200 ;
      LAYER met3 ;
        RECT 493.390 485.330 493.770 485.340 ;
        RECT 496.405 485.330 496.735 485.345 ;
        RECT 493.390 485.030 496.735 485.330 ;
        RECT 493.390 485.020 493.770 485.030 ;
        RECT 496.405 485.015 496.735 485.030 ;
        RECT 493.390 122.210 493.770 122.220 ;
        RECT 765.965 122.210 766.295 122.225 ;
        RECT 493.390 121.910 766.295 122.210 ;
        RECT 493.390 121.900 493.770 121.910 ;
        RECT 765.965 121.895 766.295 121.910 ;
      LAYER via3 ;
        RECT 493.420 485.020 493.740 485.340 ;
        RECT 493.420 121.900 493.740 122.220 ;
      LAYER met4 ;
        RECT 493.415 485.015 493.745 485.345 ;
        RECT 493.430 122.225 493.730 485.015 ;
        RECT 493.415 121.895 493.745 122.225 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.730 491.540 608.050 491.600 ;
        RECT 609.570 491.540 609.890 491.600 ;
        RECT 607.730 491.400 609.890 491.540 ;
        RECT 607.730 491.340 608.050 491.400 ;
        RECT 609.570 491.340 609.890 491.400 ;
        RECT 607.730 94.420 608.050 94.480 ;
        RECT 2221.870 94.420 2222.190 94.480 ;
        RECT 607.730 94.280 2222.190 94.420 ;
        RECT 607.730 94.220 608.050 94.280 ;
        RECT 2221.870 94.220 2222.190 94.280 ;
      LAYER via ;
        RECT 607.760 491.340 608.020 491.600 ;
        RECT 609.600 491.340 609.860 491.600 ;
        RECT 607.760 94.220 608.020 94.480 ;
        RECT 2221.900 94.220 2222.160 94.480 ;
      LAYER met2 ;
        RECT 609.390 500.000 609.670 504.000 ;
        RECT 609.430 498.680 609.570 500.000 ;
        RECT 609.430 498.540 609.800 498.680 ;
        RECT 609.660 491.630 609.800 498.540 ;
        RECT 607.760 491.310 608.020 491.630 ;
        RECT 609.600 491.310 609.860 491.630 ;
        RECT 607.820 94.510 607.960 491.310 ;
        RECT 607.760 94.190 608.020 94.510 ;
        RECT 2221.900 94.190 2222.160 94.510 ;
        RECT 2221.960 82.870 2222.100 94.190 ;
        RECT 2221.960 82.730 2225.320 82.870 ;
        RECT 2225.180 2.400 2225.320 82.730 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 608.190 472.500 608.510 472.560 ;
        RECT 610.950 472.500 611.270 472.560 ;
        RECT 608.190 472.360 611.270 472.500 ;
        RECT 608.190 472.300 608.510 472.360 ;
        RECT 610.950 472.300 611.270 472.360 ;
        RECT 608.190 100.880 608.510 100.940 ;
        RECT 2242.570 100.880 2242.890 100.940 ;
        RECT 608.190 100.740 2242.890 100.880 ;
        RECT 608.190 100.680 608.510 100.740 ;
        RECT 2242.570 100.680 2242.890 100.740 ;
      LAYER via ;
        RECT 608.220 472.300 608.480 472.560 ;
        RECT 610.980 472.300 611.240 472.560 ;
        RECT 608.220 100.680 608.480 100.940 ;
        RECT 2242.600 100.680 2242.860 100.940 ;
      LAYER met2 ;
        RECT 610.770 500.000 611.050 504.000 ;
        RECT 610.810 498.680 610.950 500.000 ;
        RECT 610.810 498.540 611.180 498.680 ;
        RECT 611.040 472.590 611.180 498.540 ;
        RECT 608.220 472.270 608.480 472.590 ;
        RECT 610.980 472.270 611.240 472.590 ;
        RECT 608.280 100.970 608.420 472.270 ;
        RECT 608.220 100.650 608.480 100.970 ;
        RECT 2242.600 100.650 2242.860 100.970 ;
        RECT 2242.660 16.050 2242.800 100.650 ;
        RECT 2242.660 15.910 2243.260 16.050 ;
        RECT 2243.120 2.400 2243.260 15.910 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.150 500.000 612.430 504.000 ;
        RECT 612.190 498.850 612.330 500.000 ;
        RECT 612.190 498.710 612.560 498.850 ;
        RECT 612.420 483.325 612.560 498.710 ;
        RECT 612.350 482.955 612.630 483.325 ;
        RECT 2256.390 100.115 2256.670 100.485 ;
        RECT 2256.460 82.870 2256.600 100.115 ;
        RECT 2256.460 82.730 2258.440 82.870 ;
        RECT 2258.300 1.770 2258.440 82.730 ;
        RECT 2260.390 1.770 2260.950 2.400 ;
        RECT 2258.300 1.630 2260.950 1.770 ;
        RECT 2260.390 -4.800 2260.950 1.630 ;
      LAYER via2 ;
        RECT 612.350 483.000 612.630 483.280 ;
        RECT 2256.390 100.160 2256.670 100.440 ;
      LAYER met3 ;
        RECT 612.325 483.290 612.655 483.305 ;
        RECT 612.990 483.290 613.370 483.300 ;
        RECT 612.325 482.990 613.370 483.290 ;
        RECT 612.325 482.975 612.655 482.990 ;
        RECT 612.990 482.980 613.370 482.990 ;
        RECT 612.990 100.450 613.370 100.460 ;
        RECT 2256.365 100.450 2256.695 100.465 ;
        RECT 612.990 100.150 2256.695 100.450 ;
        RECT 612.990 100.140 613.370 100.150 ;
        RECT 2256.365 100.135 2256.695 100.150 ;
      LAYER via3 ;
        RECT 613.020 482.980 613.340 483.300 ;
        RECT 613.020 100.140 613.340 100.460 ;
      LAYER met4 ;
        RECT 613.015 482.975 613.345 483.305 ;
        RECT 613.030 100.465 613.330 482.975 ;
        RECT 613.015 100.135 613.345 100.465 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 613.480 499.160 613.800 499.420 ;
        RECT 613.570 498.400 613.710 499.160 ;
        RECT 613.250 498.200 613.710 498.400 ;
        RECT 613.250 498.140 613.570 498.200 ;
      LAYER via ;
        RECT 613.510 499.160 613.770 499.420 ;
        RECT 613.280 498.140 613.540 498.400 ;
      LAYER met2 ;
        RECT 613.530 500.000 613.810 504.000 ;
        RECT 613.570 499.450 613.710 500.000 ;
        RECT 613.510 499.130 613.770 499.450 ;
        RECT 613.280 498.110 613.540 498.430 ;
        RECT 613.340 484.005 613.480 498.110 ;
        RECT 613.270 483.635 613.550 484.005 ;
        RECT 2277.090 121.195 2277.370 121.565 ;
        RECT 2277.160 82.870 2277.300 121.195 ;
        RECT 2277.160 82.730 2278.680 82.870 ;
        RECT 2278.540 2.400 2278.680 82.730 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
      LAYER via2 ;
        RECT 613.270 483.680 613.550 483.960 ;
        RECT 2277.090 121.240 2277.370 121.520 ;
      LAYER met3 ;
        RECT 612.070 483.970 612.450 483.980 ;
        RECT 613.245 483.970 613.575 483.985 ;
        RECT 612.070 483.670 613.575 483.970 ;
        RECT 612.070 483.660 612.450 483.670 ;
        RECT 613.245 483.655 613.575 483.670 ;
        RECT 612.070 121.530 612.450 121.540 ;
        RECT 2277.065 121.530 2277.395 121.545 ;
        RECT 612.070 121.230 2277.395 121.530 ;
        RECT 612.070 121.220 612.450 121.230 ;
        RECT 2277.065 121.215 2277.395 121.230 ;
      LAYER via3 ;
        RECT 612.100 483.660 612.420 483.980 ;
        RECT 612.100 121.220 612.420 121.540 ;
      LAYER met4 ;
        RECT 612.095 483.655 612.425 483.985 ;
        RECT 612.110 121.545 612.410 483.655 ;
        RECT 612.095 121.215 612.425 121.545 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 665.230 501.060 665.550 501.120 ;
        RECT 614.950 500.920 665.550 501.060 ;
        RECT 614.950 499.760 615.090 500.920 ;
        RECT 665.230 500.860 665.550 500.920 ;
        RECT 614.860 499.500 615.180 499.760 ;
        RECT 665.230 497.320 665.550 497.380 ;
        RECT 2290.870 497.320 2291.190 497.380 ;
        RECT 665.230 497.180 2291.190 497.320 ;
        RECT 665.230 497.120 665.550 497.180 ;
        RECT 2290.870 497.120 2291.190 497.180 ;
      LAYER via ;
        RECT 665.260 500.860 665.520 501.120 ;
        RECT 614.890 499.500 615.150 499.760 ;
        RECT 665.260 497.120 665.520 497.380 ;
        RECT 2290.900 497.120 2291.160 497.380 ;
      LAYER met2 ;
        RECT 614.910 500.000 615.190 504.000 ;
        RECT 665.260 500.830 665.520 501.150 ;
        RECT 614.950 499.790 615.090 500.000 ;
        RECT 614.890 499.470 615.150 499.790 ;
        RECT 665.320 497.410 665.460 500.830 ;
        RECT 665.260 497.090 665.520 497.410 ;
        RECT 2290.900 497.090 2291.160 497.410 ;
        RECT 2290.960 82.870 2291.100 497.090 ;
        RECT 2290.960 82.730 2296.160 82.870 ;
        RECT 2296.020 2.400 2296.160 82.730 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 616.240 500.720 616.560 500.780 ;
        RECT 616.240 500.580 646.370 500.720 ;
        RECT 616.240 500.520 616.560 500.580 ;
        RECT 646.230 500.040 646.370 500.580 ;
        RECT 666.610 500.380 666.930 500.440 ;
        RECT 647.150 500.240 666.930 500.380 ;
        RECT 647.150 500.040 647.290 500.240 ;
        RECT 666.610 500.180 666.930 500.240 ;
        RECT 646.230 499.900 647.290 500.040 ;
        RECT 666.610 496.980 666.930 497.040 ;
        RECT 2311.570 496.980 2311.890 497.040 ;
        RECT 666.610 496.840 2311.890 496.980 ;
        RECT 666.610 496.780 666.930 496.840 ;
        RECT 2311.570 496.780 2311.890 496.840 ;
      LAYER via ;
        RECT 616.270 500.520 616.530 500.780 ;
        RECT 666.640 500.180 666.900 500.440 ;
        RECT 666.640 496.780 666.900 497.040 ;
        RECT 2311.600 496.780 2311.860 497.040 ;
      LAYER met2 ;
        RECT 616.290 500.810 616.570 504.000 ;
        RECT 616.270 500.490 616.570 500.810 ;
        RECT 616.290 500.000 616.570 500.490 ;
        RECT 666.640 500.150 666.900 500.470 ;
        RECT 666.700 497.070 666.840 500.150 ;
        RECT 666.640 496.750 666.900 497.070 ;
        RECT 2311.600 496.750 2311.860 497.070 ;
        RECT 2311.660 1.770 2311.800 496.750 ;
        RECT 2313.750 1.770 2314.310 2.400 ;
        RECT 2311.660 1.630 2314.310 1.770 ;
        RECT 2313.750 -4.800 2314.310 1.630 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 617.620 499.160 617.940 499.420 ;
        RECT 614.170 497.660 614.490 497.720 ;
        RECT 617.710 497.660 617.850 499.160 ;
        RECT 614.170 497.520 617.850 497.660 ;
        RECT 614.170 497.460 614.490 497.520 ;
        RECT 614.170 86.260 614.490 86.320 ;
        RECT 2325.830 86.260 2326.150 86.320 ;
        RECT 614.170 86.120 2326.150 86.260 ;
        RECT 614.170 86.060 614.490 86.120 ;
        RECT 2325.830 86.060 2326.150 86.120 ;
      LAYER via ;
        RECT 617.650 499.160 617.910 499.420 ;
        RECT 614.200 497.460 614.460 497.720 ;
        RECT 614.200 86.060 614.460 86.320 ;
        RECT 2325.860 86.060 2326.120 86.320 ;
      LAYER met2 ;
        RECT 617.670 500.000 617.950 504.000 ;
        RECT 617.710 499.450 617.850 500.000 ;
        RECT 617.650 499.130 617.910 499.450 ;
        RECT 614.200 497.430 614.460 497.750 ;
        RECT 614.260 86.350 614.400 497.430 ;
        RECT 614.200 86.030 614.460 86.350 ;
        RECT 2325.860 86.030 2326.120 86.350 ;
        RECT 2325.920 82.870 2326.060 86.030 ;
        RECT 2325.920 82.730 2328.360 82.870 ;
        RECT 2328.220 34.570 2328.360 82.730 ;
        RECT 2328.220 34.430 2329.280 34.570 ;
        RECT 2329.140 1.770 2329.280 34.430 ;
        RECT 2331.230 1.770 2331.790 2.400 ;
        RECT 2329.140 1.630 2331.790 1.770 ;
        RECT 2331.230 -4.800 2331.790 1.630 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 615.090 472.500 615.410 472.560 ;
        RECT 619.230 472.500 619.550 472.560 ;
        RECT 615.090 472.360 619.550 472.500 ;
        RECT 615.090 472.300 615.410 472.360 ;
        RECT 619.230 472.300 619.550 472.360 ;
        RECT 615.090 128.080 615.410 128.140 ;
        RECT 2346.070 128.080 2346.390 128.140 ;
        RECT 615.090 127.940 2346.390 128.080 ;
        RECT 615.090 127.880 615.410 127.940 ;
        RECT 2346.070 127.880 2346.390 127.940 ;
      LAYER via ;
        RECT 615.120 472.300 615.380 472.560 ;
        RECT 619.260 472.300 619.520 472.560 ;
        RECT 615.120 127.880 615.380 128.140 ;
        RECT 2346.100 127.880 2346.360 128.140 ;
      LAYER met2 ;
        RECT 619.050 500.000 619.330 504.000 ;
        RECT 619.090 498.850 619.230 500.000 ;
        RECT 618.860 498.710 619.230 498.850 ;
        RECT 618.860 496.130 619.000 498.710 ;
        RECT 618.860 495.990 619.460 496.130 ;
        RECT 619.320 472.590 619.460 495.990 ;
        RECT 615.120 472.270 615.380 472.590 ;
        RECT 619.260 472.270 619.520 472.590 ;
        RECT 615.180 128.170 615.320 472.270 ;
        RECT 615.120 127.850 615.380 128.170 ;
        RECT 2346.100 127.850 2346.360 128.170 ;
        RECT 2346.160 82.870 2346.300 127.850 ;
        RECT 2346.160 82.730 2349.520 82.870 ;
        RECT 2349.380 2.400 2349.520 82.730 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.430 500.000 620.710 504.000 ;
        RECT 620.470 499.645 620.610 500.000 ;
        RECT 620.400 499.275 620.680 499.645 ;
        RECT 2367.250 128.675 2367.530 129.045 ;
        RECT 2367.320 2.400 2367.460 128.675 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
      LAYER via2 ;
        RECT 620.400 499.320 620.680 499.600 ;
        RECT 2367.250 128.720 2367.530 129.000 ;
      LAYER met3 ;
        RECT 614.830 499.610 615.210 499.620 ;
        RECT 620.375 499.610 620.705 499.625 ;
        RECT 614.830 499.310 620.705 499.610 ;
        RECT 614.830 499.300 615.210 499.310 ;
        RECT 620.375 499.295 620.705 499.310 ;
        RECT 614.830 129.010 615.210 129.020 ;
        RECT 2367.225 129.010 2367.555 129.025 ;
        RECT 614.830 128.710 2367.555 129.010 ;
        RECT 614.830 128.700 615.210 128.710 ;
        RECT 2367.225 128.695 2367.555 128.710 ;
      LAYER via3 ;
        RECT 614.860 499.300 615.180 499.620 ;
        RECT 614.860 128.700 615.180 129.020 ;
      LAYER met4 ;
        RECT 614.855 499.295 615.185 499.625 ;
        RECT 614.870 129.025 615.170 499.295 ;
        RECT 614.855 128.695 615.185 129.025 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.450 72.320 622.770 72.380 ;
        RECT 2382.410 72.320 2382.730 72.380 ;
        RECT 622.450 72.180 2382.730 72.320 ;
        RECT 622.450 72.120 622.770 72.180 ;
        RECT 2382.410 72.120 2382.730 72.180 ;
      LAYER via ;
        RECT 622.480 72.120 622.740 72.380 ;
        RECT 2382.440 72.120 2382.700 72.380 ;
      LAYER met2 ;
        RECT 621.810 500.000 622.090 504.000 ;
        RECT 621.850 498.680 621.990 500.000 ;
        RECT 621.850 498.540 622.680 498.680 ;
        RECT 622.540 72.410 622.680 498.540 ;
        RECT 622.480 72.090 622.740 72.410 ;
        RECT 2382.440 72.090 2382.700 72.410 ;
        RECT 2382.500 1.770 2382.640 72.090 ;
        RECT 2384.590 1.770 2385.150 2.400 ;
        RECT 2382.500 1.630 2385.150 1.770 ;
        RECT 2384.590 -4.800 2385.150 1.630 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.560 498.820 497.880 499.080 ;
        RECT 497.650 498.680 497.790 498.820 ;
        RECT 497.420 498.540 497.790 498.680 ;
        RECT 497.420 497.320 497.560 498.540 ;
        RECT 498.710 497.320 499.030 497.380 ;
        RECT 497.420 497.180 499.030 497.320 ;
        RECT 498.710 497.120 499.030 497.180 ;
        RECT 498.710 107.680 499.030 107.740 ;
        RECT 786.670 107.680 786.990 107.740 ;
        RECT 498.710 107.540 786.990 107.680 ;
        RECT 498.710 107.480 499.030 107.540 ;
        RECT 786.670 107.480 786.990 107.540 ;
      LAYER via ;
        RECT 497.590 498.820 497.850 499.080 ;
        RECT 498.740 497.120 499.000 497.380 ;
        RECT 498.740 107.480 499.000 107.740 ;
        RECT 786.700 107.480 786.960 107.740 ;
      LAYER met2 ;
        RECT 497.610 500.000 497.890 504.000 ;
        RECT 497.650 499.110 497.790 500.000 ;
        RECT 497.590 498.790 497.850 499.110 ;
        RECT 498.740 497.090 499.000 497.410 ;
        RECT 498.800 107.770 498.940 497.090 ;
        RECT 498.740 107.450 499.000 107.770 ;
        RECT 786.700 107.450 786.960 107.770 ;
        RECT 786.760 82.870 786.900 107.450 ;
        RECT 786.760 82.730 789.200 82.870 ;
        RECT 789.060 2.400 789.200 82.730 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 485.600 499.500 485.920 499.760 ;
        RECT 485.690 499.360 485.830 499.500 ;
        RECT 485.690 499.220 486.980 499.360 ;
        RECT 484.910 496.980 485.230 497.040 ;
        RECT 486.840 496.980 486.980 499.220 ;
        RECT 484.910 496.840 486.980 496.980 ;
        RECT 484.910 496.780 485.230 496.840 ;
        RECT 634.870 20.300 635.190 20.360 ;
        RECT 517.430 20.160 635.190 20.300 ;
        RECT 484.910 19.960 485.230 20.020 ;
        RECT 517.430 19.960 517.570 20.160 ;
        RECT 634.870 20.100 635.190 20.160 ;
        RECT 484.910 19.820 517.570 19.960 ;
        RECT 484.910 19.760 485.230 19.820 ;
      LAYER via ;
        RECT 485.630 499.500 485.890 499.760 ;
        RECT 484.940 496.780 485.200 497.040 ;
        RECT 484.940 19.760 485.200 20.020 ;
        RECT 634.900 20.100 635.160 20.360 ;
      LAYER met2 ;
        RECT 485.650 500.000 485.930 504.000 ;
        RECT 485.690 499.790 485.830 500.000 ;
        RECT 485.630 499.470 485.890 499.790 ;
        RECT 484.940 496.750 485.200 497.070 ;
        RECT 485.000 20.050 485.140 496.750 ;
        RECT 634.900 20.070 635.160 20.390 ;
        RECT 484.940 19.730 485.200 20.050 ;
        RECT 634.960 2.400 635.100 20.070 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 623.600 499.500 623.920 499.760 ;
        RECT 621.070 497.320 621.390 497.380 ;
        RECT 623.690 497.320 623.830 499.500 ;
        RECT 621.070 497.180 623.830 497.320 ;
        RECT 621.070 497.120 621.390 497.180 ;
        RECT 621.530 44.780 621.850 44.840 ;
        RECT 2408.630 44.780 2408.950 44.840 ;
        RECT 621.530 44.640 2408.950 44.780 ;
        RECT 621.530 44.580 621.850 44.640 ;
        RECT 2408.630 44.580 2408.950 44.640 ;
      LAYER via ;
        RECT 623.630 499.500 623.890 499.760 ;
        RECT 621.100 497.120 621.360 497.380 ;
        RECT 621.560 44.580 621.820 44.840 ;
        RECT 2408.660 44.580 2408.920 44.840 ;
      LAYER met2 ;
        RECT 623.650 500.000 623.930 504.000 ;
        RECT 623.690 499.790 623.830 500.000 ;
        RECT 623.630 499.470 623.890 499.790 ;
        RECT 621.100 497.090 621.360 497.410 ;
        RECT 621.160 478.450 621.300 497.090 ;
        RECT 621.160 478.310 621.760 478.450 ;
        RECT 621.620 44.870 621.760 478.310 ;
        RECT 621.560 44.550 621.820 44.870 ;
        RECT 2408.660 44.550 2408.920 44.870 ;
        RECT 2408.720 2.400 2408.860 44.550 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.990 473.520 622.310 473.580 ;
        RECT 624.290 473.520 624.610 473.580 ;
        RECT 621.990 473.380 624.610 473.520 ;
        RECT 621.990 473.320 622.310 473.380 ;
        RECT 624.290 473.320 624.610 473.380 ;
        RECT 621.990 65.520 622.310 65.580 ;
        RECT 2423.810 65.520 2424.130 65.580 ;
        RECT 621.990 65.380 2424.130 65.520 ;
        RECT 621.990 65.320 622.310 65.380 ;
        RECT 2423.810 65.320 2424.130 65.380 ;
      LAYER via ;
        RECT 622.020 473.320 622.280 473.580 ;
        RECT 624.320 473.320 624.580 473.580 ;
        RECT 622.020 65.320 622.280 65.580 ;
        RECT 2423.840 65.320 2424.100 65.580 ;
      LAYER met2 ;
        RECT 625.030 500.000 625.310 504.000 ;
        RECT 625.070 498.965 625.210 500.000 ;
        RECT 625.000 498.595 625.280 498.965 ;
        RECT 624.310 497.235 624.590 497.605 ;
        RECT 624.380 473.610 624.520 497.235 ;
        RECT 622.020 473.290 622.280 473.610 ;
        RECT 624.320 473.290 624.580 473.610 ;
        RECT 622.080 65.610 622.220 473.290 ;
        RECT 622.020 65.290 622.280 65.610 ;
        RECT 2423.840 65.290 2424.100 65.610 ;
        RECT 2423.900 1.770 2424.040 65.290 ;
        RECT 2425.990 1.770 2426.550 2.400 ;
        RECT 2423.900 1.630 2426.550 1.770 ;
        RECT 2425.990 -4.800 2426.550 1.630 ;
      LAYER via2 ;
        RECT 625.000 498.640 625.280 498.920 ;
        RECT 624.310 497.280 624.590 497.560 ;
      LAYER met3 ;
        RECT 624.975 498.615 625.305 498.945 ;
        RECT 624.285 497.570 624.615 497.585 ;
        RECT 624.990 497.570 625.290 498.615 ;
        RECT 624.285 497.270 625.290 497.570 ;
        RECT 624.285 497.255 624.615 497.270 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.410 500.000 626.690 504.000 ;
        RECT 626.450 498.680 626.590 500.000 ;
        RECT 626.450 498.540 626.820 498.680 ;
        RECT 626.680 484.005 626.820 498.540 ;
        RECT 626.610 483.635 626.890 484.005 ;
        RECT 2444.070 26.675 2444.350 27.045 ;
        RECT 2444.140 2.400 2444.280 26.675 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
      LAYER via2 ;
        RECT 626.610 483.680 626.890 483.960 ;
        RECT 2444.070 26.720 2444.350 27.000 ;
      LAYER met3 ;
        RECT 624.950 483.970 625.330 483.980 ;
        RECT 626.585 483.970 626.915 483.985 ;
        RECT 624.950 483.670 626.915 483.970 ;
        RECT 624.950 483.660 625.330 483.670 ;
        RECT 626.585 483.655 626.915 483.670 ;
        RECT 624.950 27.010 625.330 27.020 ;
        RECT 2444.045 27.010 2444.375 27.025 ;
        RECT 624.950 26.710 2444.375 27.010 ;
        RECT 624.950 26.700 625.330 26.710 ;
        RECT 2444.045 26.695 2444.375 26.710 ;
      LAYER via3 ;
        RECT 624.980 483.660 625.300 483.980 ;
        RECT 624.980 26.700 625.300 27.020 ;
      LAYER met4 ;
        RECT 624.975 483.655 625.305 483.985 ;
        RECT 624.990 27.025 625.290 483.655 ;
        RECT 624.975 26.695 625.305 27.025 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 627.740 498.820 628.060 499.080 ;
        RECT 627.830 497.040 627.970 498.820 ;
        RECT 627.830 496.840 628.290 497.040 ;
        RECT 627.970 496.780 628.290 496.840 ;
        RECT 627.970 487.120 628.290 487.180 ;
        RECT 630.270 487.120 630.590 487.180 ;
        RECT 627.970 486.980 630.590 487.120 ;
        RECT 627.970 486.920 628.290 486.980 ;
        RECT 630.270 486.920 630.590 486.980 ;
        RECT 630.270 79.460 630.590 79.520 ;
        RECT 2461.530 79.460 2461.850 79.520 ;
        RECT 630.270 79.320 2461.850 79.460 ;
        RECT 630.270 79.260 630.590 79.320 ;
        RECT 2461.530 79.260 2461.850 79.320 ;
      LAYER via ;
        RECT 627.770 498.820 628.030 499.080 ;
        RECT 628.000 496.780 628.260 497.040 ;
        RECT 628.000 486.920 628.260 487.180 ;
        RECT 630.300 486.920 630.560 487.180 ;
        RECT 630.300 79.260 630.560 79.520 ;
        RECT 2461.560 79.260 2461.820 79.520 ;
      LAYER met2 ;
        RECT 627.790 500.000 628.070 504.000 ;
        RECT 627.830 499.110 627.970 500.000 ;
        RECT 627.770 498.790 628.030 499.110 ;
        RECT 628.000 496.750 628.260 497.070 ;
        RECT 628.060 487.210 628.200 496.750 ;
        RECT 628.000 486.890 628.260 487.210 ;
        RECT 630.300 486.890 630.560 487.210 ;
        RECT 630.360 79.550 630.500 486.890 ;
        RECT 630.300 79.230 630.560 79.550 ;
        RECT 2461.560 79.230 2461.820 79.550 ;
        RECT 2461.620 2.400 2461.760 79.230 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 628.890 25.060 629.210 25.120 ;
        RECT 2479.470 25.060 2479.790 25.120 ;
        RECT 628.890 24.920 2479.790 25.060 ;
        RECT 628.890 24.860 629.210 24.920 ;
        RECT 2479.470 24.860 2479.790 24.920 ;
      LAYER via ;
        RECT 628.920 24.860 629.180 25.120 ;
        RECT 2479.500 24.860 2479.760 25.120 ;
      LAYER met2 ;
        RECT 629.170 500.000 629.450 504.000 ;
        RECT 629.210 498.340 629.350 500.000 ;
        RECT 628.980 498.200 629.350 498.340 ;
        RECT 628.980 25.150 629.120 498.200 ;
        RECT 628.920 24.830 629.180 25.150 ;
        RECT 2479.500 24.830 2479.760 25.150 ;
        RECT 2479.560 2.400 2479.700 24.830 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 629.810 33.560 630.130 33.620 ;
        RECT 2496.950 33.560 2497.270 33.620 ;
        RECT 629.810 33.420 2497.270 33.560 ;
        RECT 629.810 33.360 630.130 33.420 ;
        RECT 2496.950 33.360 2497.270 33.420 ;
      LAYER via ;
        RECT 629.840 33.360 630.100 33.620 ;
        RECT 2496.980 33.360 2497.240 33.620 ;
      LAYER met2 ;
        RECT 630.550 500.000 630.830 504.000 ;
        RECT 630.590 498.850 630.730 500.000 ;
        RECT 629.900 498.710 630.730 498.850 ;
        RECT 629.900 33.650 630.040 498.710 ;
        RECT 629.840 33.330 630.100 33.650 ;
        RECT 2496.980 33.330 2497.240 33.650 ;
        RECT 2497.040 2.400 2497.180 33.330 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 631.880 499.160 632.200 499.420 ;
        RECT 629.350 497.660 629.670 497.720 ;
        RECT 631.970 497.660 632.110 499.160 ;
        RECT 629.350 497.520 632.110 497.660 ;
        RECT 629.350 497.460 629.670 497.520 ;
        RECT 629.350 33.220 629.670 33.280 ;
        RECT 2514.890 33.220 2515.210 33.280 ;
        RECT 629.350 33.080 2515.210 33.220 ;
        RECT 629.350 33.020 629.670 33.080 ;
        RECT 2514.890 33.020 2515.210 33.080 ;
      LAYER via ;
        RECT 631.910 499.160 632.170 499.420 ;
        RECT 629.380 497.460 629.640 497.720 ;
        RECT 629.380 33.020 629.640 33.280 ;
        RECT 2514.920 33.020 2515.180 33.280 ;
      LAYER met2 ;
        RECT 631.930 500.000 632.210 504.000 ;
        RECT 631.970 499.450 632.110 500.000 ;
        RECT 631.910 499.130 632.170 499.450 ;
        RECT 629.380 497.430 629.640 497.750 ;
        RECT 629.440 33.310 629.580 497.430 ;
        RECT 629.380 32.990 629.640 33.310 ;
        RECT 2514.920 32.990 2515.180 33.310 ;
        RECT 2514.980 2.400 2515.120 32.990 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.310 500.000 633.590 504.000 ;
        RECT 633.350 498.850 633.490 500.000 ;
        RECT 633.350 498.710 633.720 498.850 ;
        RECT 633.580 483.325 633.720 498.710 ;
        RECT 633.510 482.955 633.790 483.325 ;
        RECT 2532.850 79.035 2533.130 79.405 ;
        RECT 2532.920 16.730 2533.060 79.035 ;
        RECT 2532.460 16.590 2533.060 16.730 ;
        RECT 2532.460 2.400 2532.600 16.590 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
      LAYER via2 ;
        RECT 633.510 483.000 633.790 483.280 ;
        RECT 2532.850 79.080 2533.130 79.360 ;
      LAYER met3 ;
        RECT 633.485 483.300 633.815 483.305 ;
        RECT 633.230 483.290 633.815 483.300 ;
        RECT 633.030 482.990 633.815 483.290 ;
        RECT 633.230 482.980 633.815 482.990 ;
        RECT 633.485 482.975 633.815 482.980 ;
        RECT 633.230 79.370 633.610 79.380 ;
        RECT 2532.825 79.370 2533.155 79.385 ;
        RECT 633.230 79.070 2533.155 79.370 ;
        RECT 633.230 79.060 633.610 79.070 ;
        RECT 2532.825 79.055 2533.155 79.070 ;
      LAYER via3 ;
        RECT 633.260 482.980 633.580 483.300 ;
        RECT 633.260 79.060 633.580 79.380 ;
      LAYER met4 ;
        RECT 633.255 482.975 633.585 483.305 ;
        RECT 633.270 79.385 633.570 482.975 ;
        RECT 633.255 79.055 633.585 79.385 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.410 498.000 634.730 498.060 ;
        RECT 635.330 498.000 635.650 498.060 ;
        RECT 634.410 497.860 635.650 498.000 ;
        RECT 634.410 497.800 634.730 497.860 ;
        RECT 635.330 497.800 635.650 497.860 ;
        RECT 635.330 100.540 635.650 100.600 ;
        RECT 2546.170 100.540 2546.490 100.600 ;
        RECT 635.330 100.400 2546.490 100.540 ;
        RECT 635.330 100.340 635.650 100.400 ;
        RECT 2546.170 100.340 2546.490 100.400 ;
      LAYER via ;
        RECT 634.440 497.800 634.700 498.060 ;
        RECT 635.360 497.800 635.620 498.060 ;
        RECT 635.360 100.340 635.620 100.600 ;
        RECT 2546.200 100.340 2546.460 100.600 ;
      LAYER met2 ;
        RECT 634.690 500.000 634.970 504.000 ;
        RECT 634.730 499.020 634.870 500.000 ;
        RECT 634.500 498.880 634.870 499.020 ;
        RECT 634.500 498.090 634.640 498.880 ;
        RECT 634.440 497.770 634.700 498.090 ;
        RECT 635.360 497.770 635.620 498.090 ;
        RECT 635.420 100.630 635.560 497.770 ;
        RECT 635.360 100.310 635.620 100.630 ;
        RECT 2546.200 100.310 2546.460 100.630 ;
        RECT 2546.260 82.870 2546.400 100.310 ;
        RECT 2546.260 82.730 2548.240 82.870 ;
        RECT 2548.100 1.770 2548.240 82.730 ;
        RECT 2550.190 1.770 2550.750 2.400 ;
        RECT 2548.100 1.630 2550.750 1.770 ;
        RECT 2550.190 -4.800 2550.750 1.630 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 636.020 499.500 636.340 499.760 ;
        RECT 636.110 499.080 636.250 499.500 ;
        RECT 635.790 498.880 636.250 499.080 ;
        RECT 635.790 498.820 636.110 498.880 ;
        RECT 635.790 107.340 636.110 107.400 ;
        RECT 2566.870 107.340 2567.190 107.400 ;
        RECT 635.790 107.200 2567.190 107.340 ;
        RECT 635.790 107.140 636.110 107.200 ;
        RECT 2566.870 107.140 2567.190 107.200 ;
      LAYER via ;
        RECT 636.050 499.500 636.310 499.760 ;
        RECT 635.820 498.820 636.080 499.080 ;
        RECT 635.820 107.140 636.080 107.400 ;
        RECT 2566.900 107.140 2567.160 107.400 ;
      LAYER met2 ;
        RECT 636.070 500.000 636.350 504.000 ;
        RECT 636.110 499.790 636.250 500.000 ;
        RECT 636.050 499.470 636.310 499.790 ;
        RECT 635.820 498.790 636.080 499.110 ;
        RECT 635.880 107.430 636.020 498.790 ;
        RECT 635.820 107.110 636.080 107.430 ;
        RECT 2566.900 107.110 2567.160 107.430 ;
        RECT 2566.960 1.770 2567.100 107.110 ;
        RECT 2567.670 1.770 2568.230 2.400 ;
        RECT 2566.960 1.630 2568.230 1.770 ;
        RECT 2567.670 -4.800 2568.230 1.630 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.330 472.840 497.650 472.900 ;
        RECT 499.630 472.840 499.950 472.900 ;
        RECT 497.330 472.700 499.950 472.840 ;
        RECT 497.330 472.640 497.650 472.700 ;
        RECT 499.630 472.640 499.950 472.700 ;
        RECT 497.330 25.400 497.650 25.460 ;
        RECT 812.430 25.400 812.750 25.460 ;
        RECT 497.330 25.260 812.750 25.400 ;
        RECT 497.330 25.200 497.650 25.260 ;
        RECT 812.430 25.200 812.750 25.260 ;
      LAYER via ;
        RECT 497.360 472.640 497.620 472.900 ;
        RECT 499.660 472.640 499.920 472.900 ;
        RECT 497.360 25.200 497.620 25.460 ;
        RECT 812.460 25.200 812.720 25.460 ;
      LAYER met2 ;
        RECT 499.450 500.000 499.730 504.000 ;
        RECT 499.490 498.340 499.630 500.000 ;
        RECT 499.490 498.200 499.860 498.340 ;
        RECT 499.720 472.930 499.860 498.200 ;
        RECT 497.360 472.610 497.620 472.930 ;
        RECT 499.660 472.610 499.920 472.930 ;
        RECT 497.420 25.490 497.560 472.610 ;
        RECT 497.360 25.170 497.620 25.490 ;
        RECT 812.460 25.170 812.720 25.490 ;
        RECT 812.520 2.400 812.660 25.170 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 637.400 499.500 637.720 499.760 ;
        RECT 637.490 499.080 637.630 499.500 ;
        RECT 637.170 498.880 637.630 499.080 ;
        RECT 637.170 498.820 637.490 498.880 ;
        RECT 636.250 107.000 636.570 107.060 ;
        RECT 2580.670 107.000 2580.990 107.060 ;
        RECT 636.250 106.860 2580.990 107.000 ;
        RECT 636.250 106.800 636.570 106.860 ;
        RECT 2580.670 106.800 2580.990 106.860 ;
      LAYER via ;
        RECT 637.430 499.500 637.690 499.760 ;
        RECT 637.200 498.820 637.460 499.080 ;
        RECT 636.280 106.800 636.540 107.060 ;
        RECT 2580.700 106.800 2580.960 107.060 ;
      LAYER met2 ;
        RECT 637.450 500.000 637.730 504.000 ;
        RECT 637.490 499.790 637.630 500.000 ;
        RECT 637.430 499.470 637.690 499.790 ;
        RECT 637.200 499.020 637.460 499.110 ;
        RECT 636.800 498.880 637.460 499.020 ;
        RECT 636.800 473.010 636.940 498.880 ;
        RECT 637.200 498.790 637.460 498.880 ;
        RECT 636.340 472.870 636.940 473.010 ;
        RECT 636.340 107.090 636.480 472.870 ;
        RECT 636.280 106.770 636.540 107.090 ;
        RECT 2580.700 106.770 2580.960 107.090 ;
        RECT 2580.760 82.870 2580.900 106.770 ;
        RECT 2580.760 82.730 2585.960 82.870 ;
        RECT 2585.820 2.400 2585.960 82.730 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 638.780 499.500 639.100 499.760 ;
        RECT 637.170 497.660 637.490 497.720 ;
        RECT 638.870 497.660 639.010 499.500 ;
        RECT 637.170 497.520 639.010 497.660 ;
        RECT 637.170 497.460 637.490 497.520 ;
        RECT 636.710 114.140 637.030 114.200 ;
        RECT 2601.370 114.140 2601.690 114.200 ;
        RECT 636.710 114.000 2601.690 114.140 ;
        RECT 636.710 113.940 637.030 114.000 ;
        RECT 2601.370 113.940 2601.690 114.000 ;
      LAYER via ;
        RECT 638.810 499.500 639.070 499.760 ;
        RECT 637.200 497.460 637.460 497.720 ;
        RECT 636.740 113.940 637.000 114.200 ;
        RECT 2601.400 113.940 2601.660 114.200 ;
      LAYER met2 ;
        RECT 638.830 500.000 639.110 504.000 ;
        RECT 638.870 499.790 639.010 500.000 ;
        RECT 638.810 499.470 639.070 499.790 ;
        RECT 637.200 497.430 637.460 497.750 ;
        RECT 637.260 472.330 637.400 497.430 ;
        RECT 636.800 472.190 637.400 472.330 ;
        RECT 636.800 114.230 636.940 472.190 ;
        RECT 636.740 113.910 637.000 114.230 ;
        RECT 2601.400 113.910 2601.660 114.230 ;
        RECT 2601.460 1.770 2601.600 113.910 ;
        RECT 2603.550 1.770 2604.110 2.400 ;
        RECT 2601.460 1.630 2604.110 1.770 ;
        RECT 2603.550 -4.800 2604.110 1.630 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.210 500.000 640.490 504.000 ;
        RECT 640.250 499.815 640.390 500.000 ;
        RECT 640.180 499.445 640.460 499.815 ;
        RECT 2615.190 127.995 2615.470 128.365 ;
        RECT 2615.260 82.870 2615.400 127.995 ;
        RECT 2615.260 82.730 2619.080 82.870 ;
        RECT 2618.940 1.770 2619.080 82.730 ;
        RECT 2621.030 1.770 2621.590 2.400 ;
        RECT 2618.940 1.630 2621.590 1.770 ;
        RECT 2621.030 -4.800 2621.590 1.630 ;
      LAYER via2 ;
        RECT 640.180 499.490 640.460 499.770 ;
        RECT 2615.190 128.040 2615.470 128.320 ;
      LAYER met3 ;
        RECT 640.155 499.780 640.485 499.795 ;
        RECT 639.940 499.465 640.485 499.780 ;
        RECT 636.910 498.250 637.290 498.260 ;
        RECT 639.940 498.250 640.240 499.465 ;
        RECT 636.910 497.950 640.240 498.250 ;
        RECT 636.910 497.940 637.290 497.950 ;
        RECT 636.910 128.330 637.290 128.340 ;
        RECT 2615.165 128.330 2615.495 128.345 ;
        RECT 636.910 128.030 2615.495 128.330 ;
        RECT 636.910 128.020 637.290 128.030 ;
        RECT 2615.165 128.015 2615.495 128.030 ;
      LAYER via3 ;
        RECT 636.940 497.940 637.260 498.260 ;
        RECT 636.940 128.020 637.260 128.340 ;
      LAYER met4 ;
        RECT 636.935 497.935 637.265 498.265 ;
        RECT 636.950 128.345 637.250 497.935 ;
        RECT 636.935 128.015 637.265 128.345 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 641.770 488.480 642.090 488.540 ;
        RECT 643.150 488.480 643.470 488.540 ;
        RECT 641.770 488.340 643.470 488.480 ;
        RECT 641.770 488.280 642.090 488.340 ;
        RECT 643.150 488.280 643.470 488.340 ;
        RECT 643.150 32.880 643.470 32.940 ;
        RECT 2639.090 32.880 2639.410 32.940 ;
        RECT 643.150 32.740 2639.410 32.880 ;
        RECT 643.150 32.680 643.470 32.740 ;
        RECT 2639.090 32.680 2639.410 32.740 ;
      LAYER via ;
        RECT 641.800 488.280 642.060 488.540 ;
        RECT 643.180 488.280 643.440 488.540 ;
        RECT 643.180 32.680 643.440 32.940 ;
        RECT 2639.120 32.680 2639.380 32.940 ;
      LAYER met2 ;
        RECT 641.590 500.000 641.870 504.000 ;
        RECT 641.630 498.680 641.770 500.000 ;
        RECT 641.630 498.540 642.000 498.680 ;
        RECT 641.860 488.570 642.000 498.540 ;
        RECT 641.800 488.250 642.060 488.570 ;
        RECT 643.180 488.250 643.440 488.570 ;
        RECT 643.240 32.970 643.380 488.250 ;
        RECT 643.180 32.650 643.440 32.970 ;
        RECT 2639.120 32.650 2639.380 32.970 ;
        RECT 2639.180 2.400 2639.320 32.650 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 643.610 473.520 643.930 473.580 ;
        RECT 643.610 473.380 644.760 473.520 ;
        RECT 643.610 473.320 643.930 473.380 ;
        RECT 644.620 472.560 644.760 473.380 ;
        RECT 644.530 472.300 644.850 472.560 ;
        RECT 644.530 113.800 644.850 113.860 ;
        RECT 2657.030 113.800 2657.350 113.860 ;
        RECT 644.530 113.660 2657.350 113.800 ;
        RECT 644.530 113.600 644.850 113.660 ;
        RECT 2657.030 113.600 2657.350 113.660 ;
      LAYER via ;
        RECT 643.640 473.320 643.900 473.580 ;
        RECT 644.560 472.300 644.820 472.560 ;
        RECT 644.560 113.600 644.820 113.860 ;
        RECT 2657.060 113.600 2657.320 113.860 ;
      LAYER met2 ;
        RECT 642.970 500.000 643.250 504.000 ;
        RECT 643.010 499.815 643.150 500.000 ;
        RECT 642.940 499.445 643.220 499.815 ;
        RECT 642.940 498.595 643.220 498.965 ;
        RECT 643.010 498.340 643.150 498.595 ;
        RECT 643.010 498.200 643.380 498.340 ;
        RECT 643.240 489.330 643.380 498.200 ;
        RECT 643.240 489.190 643.840 489.330 ;
        RECT 643.700 473.610 643.840 489.190 ;
        RECT 643.640 473.290 643.900 473.610 ;
        RECT 644.560 472.270 644.820 472.590 ;
        RECT 644.620 113.890 644.760 472.270 ;
        RECT 644.560 113.570 644.820 113.890 ;
        RECT 2657.060 113.570 2657.320 113.890 ;
        RECT 2657.120 16.730 2657.260 113.570 ;
        RECT 2656.660 16.590 2657.260 16.730 ;
        RECT 2656.660 2.400 2656.800 16.590 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
      LAYER via2 ;
        RECT 642.940 499.490 643.220 499.770 ;
        RECT 642.940 498.640 643.220 498.920 ;
      LAYER met3 ;
        RECT 642.915 499.780 643.245 499.795 ;
        RECT 642.700 499.465 643.245 499.780 ;
        RECT 642.700 498.945 643.000 499.465 ;
        RECT 642.700 498.630 643.245 498.945 ;
        RECT 642.915 498.615 643.245 498.630 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 641.770 32.200 642.090 32.260 ;
        RECT 2674.510 32.200 2674.830 32.260 ;
        RECT 641.770 32.060 2674.830 32.200 ;
        RECT 641.770 32.000 642.090 32.060 ;
        RECT 2674.510 32.000 2674.830 32.060 ;
      LAYER via ;
        RECT 641.800 32.000 642.060 32.260 ;
        RECT 2674.540 32.000 2674.800 32.260 ;
      LAYER met2 ;
        RECT 644.350 500.000 644.630 504.000 ;
        RECT 644.390 499.815 644.530 500.000 ;
        RECT 644.320 499.445 644.600 499.815 ;
        RECT 642.250 497.915 642.530 498.285 ;
        RECT 642.320 487.970 642.460 497.915 ;
        RECT 641.860 487.830 642.460 487.970 ;
        RECT 641.860 32.290 642.000 487.830 ;
        RECT 641.800 31.970 642.060 32.290 ;
        RECT 2674.540 31.970 2674.800 32.290 ;
        RECT 2674.600 2.400 2674.740 31.970 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
      LAYER via2 ;
        RECT 644.320 499.490 644.600 499.770 ;
        RECT 642.250 497.960 642.530 498.240 ;
      LAYER met3 ;
        RECT 644.295 499.465 644.625 499.795 ;
        RECT 642.225 498.250 642.555 498.265 ;
        RECT 644.310 498.250 644.610 499.465 ;
        RECT 642.225 497.950 644.610 498.250 ;
        RECT 642.225 497.935 642.555 497.950 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 644.070 472.160 644.390 472.220 ;
        RECT 645.910 472.160 646.230 472.220 ;
        RECT 644.070 472.020 646.230 472.160 ;
        RECT 644.070 471.960 644.390 472.020 ;
        RECT 645.910 471.960 646.230 472.020 ;
        RECT 644.070 40.020 644.390 40.080 ;
        RECT 2691.990 40.020 2692.310 40.080 ;
        RECT 644.070 39.880 2692.310 40.020 ;
        RECT 644.070 39.820 644.390 39.880 ;
        RECT 2691.990 39.820 2692.310 39.880 ;
      LAYER via ;
        RECT 644.100 471.960 644.360 472.220 ;
        RECT 645.940 471.960 646.200 472.220 ;
        RECT 644.100 39.820 644.360 40.080 ;
        RECT 2692.020 39.820 2692.280 40.080 ;
      LAYER met2 ;
        RECT 645.730 500.000 646.010 504.000 ;
        RECT 645.770 498.340 645.910 500.000 ;
        RECT 645.770 498.200 646.140 498.340 ;
        RECT 646.000 472.250 646.140 498.200 ;
        RECT 644.100 471.930 644.360 472.250 ;
        RECT 645.940 471.930 646.200 472.250 ;
        RECT 644.160 40.110 644.300 471.930 ;
        RECT 644.100 39.790 644.360 40.110 ;
        RECT 2692.020 39.790 2692.280 40.110 ;
        RECT 2692.080 2.400 2692.220 39.790 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 647.060 498.820 647.380 499.080 ;
        RECT 647.150 498.060 647.290 498.820 ;
        RECT 646.830 497.860 647.290 498.060 ;
        RECT 646.830 497.800 647.150 497.860 ;
      LAYER via ;
        RECT 647.090 498.820 647.350 499.080 ;
        RECT 646.860 497.800 647.120 498.060 ;
      LAYER met2 ;
        RECT 647.110 500.000 647.390 504.000 ;
        RECT 647.150 499.110 647.290 500.000 ;
        RECT 647.090 498.790 647.350 499.110 ;
        RECT 646.860 497.770 647.120 498.090 ;
        RECT 646.920 490.125 647.060 497.770 ;
        RECT 646.850 489.755 647.130 490.125 ;
        RECT 2704.890 127.315 2705.170 127.685 ;
        RECT 2704.960 82.870 2705.100 127.315 ;
        RECT 2704.960 82.730 2710.160 82.870 ;
        RECT 2710.020 2.400 2710.160 82.730 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
      LAYER via2 ;
        RECT 646.850 489.800 647.130 490.080 ;
        RECT 2704.890 127.360 2705.170 127.640 ;
      LAYER met3 ;
        RECT 646.825 490.100 647.155 490.105 ;
        RECT 646.825 490.090 647.410 490.100 ;
        RECT 646.825 489.790 647.610 490.090 ;
        RECT 646.825 489.780 647.410 489.790 ;
        RECT 646.825 489.775 647.155 489.780 ;
        RECT 647.030 127.650 647.410 127.660 ;
        RECT 2704.865 127.650 2705.195 127.665 ;
        RECT 647.030 127.350 2705.195 127.650 ;
        RECT 647.030 127.340 647.410 127.350 ;
        RECT 2704.865 127.335 2705.195 127.350 ;
      LAYER via3 ;
        RECT 647.060 489.780 647.380 490.100 ;
        RECT 647.060 127.340 647.380 127.660 ;
      LAYER met4 ;
        RECT 647.055 489.775 647.385 490.105 ;
        RECT 647.070 127.665 647.370 489.775 ;
        RECT 647.055 127.335 647.385 127.665 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 650.050 120.940 650.370 121.000 ;
        RECT 2725.570 120.940 2725.890 121.000 ;
        RECT 650.050 120.800 2725.890 120.940 ;
        RECT 650.050 120.740 650.370 120.800 ;
        RECT 2725.570 120.740 2725.890 120.800 ;
      LAYER via ;
        RECT 650.080 120.740 650.340 121.000 ;
        RECT 2725.600 120.740 2725.860 121.000 ;
      LAYER met2 ;
        RECT 648.490 500.000 648.770 504.000 ;
        RECT 648.530 498.680 648.670 500.000 ;
        RECT 648.530 498.540 649.360 498.680 ;
        RECT 649.220 474.370 649.360 498.540 ;
        RECT 649.220 474.230 650.280 474.370 ;
        RECT 650.140 121.030 650.280 474.230 ;
        RECT 650.080 120.710 650.340 121.030 ;
        RECT 2725.600 120.710 2725.860 121.030 ;
        RECT 2725.660 82.870 2725.800 120.710 ;
        RECT 2725.660 82.730 2727.640 82.870 ;
        RECT 2727.500 2.400 2727.640 82.730 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 649.820 499.360 650.140 499.420 ;
        RECT 649.680 499.160 650.140 499.360 ;
        RECT 649.680 498.740 649.820 499.160 ;
        RECT 649.590 498.480 649.910 498.740 ;
        RECT 650.510 120.600 650.830 120.660 ;
        RECT 2739.830 120.600 2740.150 120.660 ;
        RECT 650.510 120.460 2740.150 120.600 ;
        RECT 650.510 120.400 650.830 120.460 ;
        RECT 2739.830 120.400 2740.150 120.460 ;
      LAYER via ;
        RECT 649.850 499.160 650.110 499.420 ;
        RECT 649.620 498.480 649.880 498.740 ;
        RECT 650.540 120.400 650.800 120.660 ;
        RECT 2739.860 120.400 2740.120 120.660 ;
      LAYER met2 ;
        RECT 649.870 500.000 650.150 504.000 ;
        RECT 649.910 499.450 650.050 500.000 ;
        RECT 649.850 499.130 650.110 499.450 ;
        RECT 649.610 498.595 649.890 498.965 ;
        RECT 649.620 498.450 649.880 498.595 ;
        RECT 650.530 497.915 650.810 498.285 ;
        RECT 650.600 120.690 650.740 497.915 ;
        RECT 650.540 120.370 650.800 120.690 ;
        RECT 2739.860 120.370 2740.120 120.690 ;
        RECT 2739.920 82.870 2740.060 120.370 ;
        RECT 2739.920 82.730 2743.280 82.870 ;
        RECT 2743.140 1.770 2743.280 82.730 ;
        RECT 2745.230 1.770 2745.790 2.400 ;
        RECT 2743.140 1.630 2745.790 1.770 ;
        RECT 2745.230 -4.800 2745.790 1.630 ;
      LAYER via2 ;
        RECT 649.610 498.640 649.890 498.920 ;
        RECT 650.530 497.960 650.810 498.240 ;
      LAYER met3 ;
        RECT 649.585 498.930 649.915 498.945 ;
        RECT 649.585 498.630 650.820 498.930 ;
        RECT 649.585 498.615 649.915 498.630 ;
        RECT 650.520 498.265 650.820 498.630 ;
        RECT 650.505 497.935 650.835 498.265 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 500.780 499.160 501.100 499.420 ;
        RECT 499.170 497.660 499.490 497.720 ;
        RECT 500.870 497.660 501.010 499.160 ;
        RECT 499.170 497.520 501.010 497.660 ;
        RECT 499.170 497.460 499.490 497.520 ;
        RECT 499.170 122.980 499.490 123.040 ;
        RECT 828.070 122.980 828.390 123.040 ;
        RECT 499.170 122.840 828.390 122.980 ;
        RECT 499.170 122.780 499.490 122.840 ;
        RECT 828.070 122.780 828.390 122.840 ;
      LAYER via ;
        RECT 500.810 499.160 501.070 499.420 ;
        RECT 499.200 497.460 499.460 497.720 ;
        RECT 499.200 122.780 499.460 123.040 ;
        RECT 828.100 122.780 828.360 123.040 ;
      LAYER met2 ;
        RECT 500.830 500.000 501.110 504.000 ;
        RECT 500.870 499.450 501.010 500.000 ;
        RECT 500.810 499.130 501.070 499.450 ;
        RECT 499.200 497.430 499.460 497.750 ;
        RECT 499.260 123.070 499.400 497.430 ;
        RECT 499.200 122.750 499.460 123.070 ;
        RECT 828.100 122.750 828.360 123.070 ;
        RECT 828.160 82.870 828.300 122.750 ;
        RECT 828.160 82.730 830.600 82.870 ;
        RECT 830.460 2.400 830.600 82.730 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 651.200 499.500 651.520 499.760 ;
        RECT 651.290 498.680 651.430 499.500 ;
        RECT 651.290 498.540 652.120 498.680 ;
        RECT 648.670 497.660 648.990 497.720 ;
        RECT 651.980 497.660 652.120 498.540 ;
        RECT 648.670 497.520 652.120 497.660 ;
        RECT 648.670 497.460 648.990 497.520 ;
        RECT 649.130 31.180 649.450 31.240 ;
        RECT 2763.290 31.180 2763.610 31.240 ;
        RECT 649.130 31.040 2763.610 31.180 ;
        RECT 649.130 30.980 649.450 31.040 ;
        RECT 2763.290 30.980 2763.610 31.040 ;
      LAYER via ;
        RECT 651.230 499.500 651.490 499.760 ;
        RECT 648.700 497.460 648.960 497.720 ;
        RECT 649.160 30.980 649.420 31.240 ;
        RECT 2763.320 30.980 2763.580 31.240 ;
      LAYER met2 ;
        RECT 651.250 500.000 651.530 504.000 ;
        RECT 651.290 499.790 651.430 500.000 ;
        RECT 651.230 499.470 651.490 499.790 ;
        RECT 648.700 497.430 648.960 497.750 ;
        RECT 648.760 473.690 648.900 497.430 ;
        RECT 648.760 473.550 649.360 473.690 ;
        RECT 649.220 31.270 649.360 473.550 ;
        RECT 649.160 30.950 649.420 31.270 ;
        RECT 2763.320 30.950 2763.580 31.270 ;
        RECT 2763.380 2.400 2763.520 30.950 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 650.970 472.160 651.290 472.220 ;
        RECT 653.270 472.160 653.590 472.220 ;
        RECT 650.970 472.020 653.590 472.160 ;
        RECT 650.970 471.960 651.290 472.020 ;
        RECT 653.270 471.960 653.590 472.020 ;
        RECT 650.970 127.740 651.290 127.800 ;
        RECT 2781.230 127.740 2781.550 127.800 ;
        RECT 650.970 127.600 2781.550 127.740 ;
        RECT 650.970 127.540 651.290 127.600 ;
        RECT 2781.230 127.540 2781.550 127.600 ;
      LAYER via ;
        RECT 651.000 471.960 651.260 472.220 ;
        RECT 653.300 471.960 653.560 472.220 ;
        RECT 651.000 127.540 651.260 127.800 ;
        RECT 2781.260 127.540 2781.520 127.800 ;
      LAYER met2 ;
        RECT 652.630 500.000 652.910 504.000 ;
        RECT 652.670 499.815 652.810 500.000 ;
        RECT 652.600 499.445 652.880 499.815 ;
        RECT 652.830 497.915 653.110 498.285 ;
        RECT 652.900 488.140 653.040 497.915 ;
        RECT 652.900 488.000 653.500 488.140 ;
        RECT 653.360 472.250 653.500 488.000 ;
        RECT 651.000 471.930 651.260 472.250 ;
        RECT 653.300 471.930 653.560 472.250 ;
        RECT 651.060 127.830 651.200 471.930 ;
        RECT 651.000 127.510 651.260 127.830 ;
        RECT 2781.260 127.510 2781.520 127.830 ;
        RECT 2781.320 16.730 2781.460 127.510 ;
        RECT 2780.860 16.590 2781.460 16.730 ;
        RECT 2780.860 2.400 2781.000 16.590 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
      LAYER via2 ;
        RECT 652.600 499.490 652.880 499.770 ;
        RECT 652.830 497.960 653.110 498.240 ;
      LAYER met3 ;
        RECT 652.575 499.465 652.905 499.795 ;
        RECT 652.590 498.265 652.890 499.465 ;
        RECT 652.590 497.950 653.135 498.265 ;
        RECT 652.805 497.935 653.135 497.950 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 653.960 498.820 654.280 499.080 ;
        RECT 654.050 498.400 654.190 498.820 ;
        RECT 653.730 498.200 654.190 498.400 ;
        RECT 653.730 498.140 654.050 498.200 ;
      LAYER via ;
        RECT 653.990 498.820 654.250 499.080 ;
        RECT 653.760 498.140 654.020 498.400 ;
      LAYER met2 ;
        RECT 654.010 500.000 654.290 504.000 ;
        RECT 654.050 499.110 654.190 500.000 ;
        RECT 653.990 498.790 654.250 499.110 ;
        RECT 653.760 498.110 654.020 498.430 ;
        RECT 653.820 487.405 653.960 498.110 ;
        RECT 653.750 487.035 654.030 487.405 ;
        RECT 2794.590 134.115 2794.870 134.485 ;
        RECT 2794.660 82.870 2794.800 134.115 ;
        RECT 2794.660 82.730 2796.640 82.870 ;
        RECT 2796.500 1.770 2796.640 82.730 ;
        RECT 2798.590 1.770 2799.150 2.400 ;
        RECT 2796.500 1.630 2799.150 1.770 ;
        RECT 2798.590 -4.800 2799.150 1.630 ;
      LAYER via2 ;
        RECT 653.750 487.080 654.030 487.360 ;
        RECT 2794.590 134.160 2794.870 134.440 ;
      LAYER met3 ;
        RECT 652.550 487.370 652.930 487.380 ;
        RECT 653.725 487.370 654.055 487.385 ;
        RECT 652.550 487.070 654.055 487.370 ;
        RECT 652.550 487.060 652.930 487.070 ;
        RECT 653.725 487.055 654.055 487.070 ;
        RECT 652.550 134.450 652.930 134.460 ;
        RECT 2794.565 134.450 2794.895 134.465 ;
        RECT 652.550 134.150 2794.895 134.450 ;
        RECT 652.550 134.140 652.930 134.150 ;
        RECT 2794.565 134.135 2794.895 134.150 ;
      LAYER via3 ;
        RECT 652.580 487.060 652.900 487.380 ;
        RECT 652.580 134.140 652.900 134.460 ;
      LAYER met4 ;
        RECT 652.575 487.055 652.905 487.385 ;
        RECT 652.590 134.465 652.890 487.055 ;
        RECT 652.575 134.135 652.905 134.465 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 664.770 486.440 665.090 486.500 ;
        RECT 2815.270 486.440 2815.590 486.500 ;
        RECT 664.770 486.300 2815.590 486.440 ;
        RECT 664.770 486.240 665.090 486.300 ;
        RECT 2815.270 486.240 2815.590 486.300 ;
      LAYER via ;
        RECT 664.800 486.240 665.060 486.500 ;
        RECT 2815.300 486.240 2815.560 486.500 ;
      LAYER met2 ;
        RECT 655.390 500.000 655.670 504.000 ;
        RECT 655.430 499.645 655.570 500.000 ;
        RECT 664.790 499.955 665.070 500.325 ;
        RECT 655.360 499.275 655.640 499.645 ;
        RECT 664.860 486.530 665.000 499.955 ;
        RECT 664.800 486.210 665.060 486.530 ;
        RECT 2815.300 486.210 2815.560 486.530 ;
        RECT 2815.360 1.770 2815.500 486.210 ;
        RECT 2816.070 1.770 2816.630 2.400 ;
        RECT 2815.360 1.630 2816.630 1.770 ;
        RECT 2816.070 -4.800 2816.630 1.630 ;
      LAYER via2 ;
        RECT 664.790 500.000 665.070 500.280 ;
        RECT 655.360 499.320 655.640 499.600 ;
      LAYER met3 ;
        RECT 664.765 500.290 665.095 500.305 ;
        RECT 657.190 499.990 665.095 500.290 ;
        RECT 655.335 499.610 655.665 499.625 ;
        RECT 657.190 499.610 657.490 499.990 ;
        RECT 664.765 499.975 665.095 499.990 ;
        RECT 655.335 499.310 657.490 499.610 ;
        RECT 655.335 499.295 655.665 499.310 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.720 499.500 657.040 499.760 ;
        RECT 656.810 499.360 656.950 499.500 ;
        RECT 656.810 499.220 657.180 499.360 ;
        RECT 655.570 498.000 655.890 498.060 ;
        RECT 657.040 498.000 657.180 499.220 ;
        RECT 655.570 497.860 657.180 498.000 ;
        RECT 655.570 497.800 655.890 497.860 ;
        RECT 655.570 30.840 655.890 30.900 ;
        RECT 2834.130 30.840 2834.450 30.900 ;
        RECT 655.570 30.700 2834.450 30.840 ;
        RECT 655.570 30.640 655.890 30.700 ;
        RECT 2834.130 30.640 2834.450 30.700 ;
      LAYER via ;
        RECT 656.750 499.500 657.010 499.760 ;
        RECT 655.600 497.800 655.860 498.060 ;
        RECT 655.600 30.640 655.860 30.900 ;
        RECT 2834.160 30.640 2834.420 30.900 ;
      LAYER met2 ;
        RECT 656.770 500.000 657.050 504.000 ;
        RECT 656.810 499.790 656.950 500.000 ;
        RECT 656.750 499.470 657.010 499.790 ;
        RECT 655.600 497.770 655.860 498.090 ;
        RECT 655.660 30.930 655.800 497.770 ;
        RECT 655.600 30.610 655.860 30.930 ;
        RECT 2834.160 30.610 2834.420 30.930 ;
        RECT 2834.220 2.400 2834.360 30.610 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.490 478.280 656.810 478.340 ;
        RECT 657.410 478.280 657.730 478.340 ;
        RECT 656.490 478.140 657.730 478.280 ;
        RECT 656.490 478.080 656.810 478.140 ;
        RECT 657.410 478.080 657.730 478.140 ;
        RECT 656.490 38.660 656.810 38.720 ;
        RECT 2851.610 38.660 2851.930 38.720 ;
        RECT 656.490 38.520 2851.930 38.660 ;
        RECT 656.490 38.460 656.810 38.520 ;
        RECT 2851.610 38.460 2851.930 38.520 ;
      LAYER via ;
        RECT 656.520 478.080 656.780 478.340 ;
        RECT 657.440 478.080 657.700 478.340 ;
        RECT 656.520 38.460 656.780 38.720 ;
        RECT 2851.640 38.460 2851.900 38.720 ;
      LAYER met2 ;
        RECT 658.150 500.000 658.430 504.000 ;
        RECT 658.190 499.475 658.330 500.000 ;
        RECT 658.120 499.105 658.400 499.475 ;
        RECT 657.430 497.235 657.710 497.605 ;
        RECT 657.500 478.370 657.640 497.235 ;
        RECT 656.520 478.050 656.780 478.370 ;
        RECT 657.440 478.050 657.700 478.370 ;
        RECT 656.580 38.750 656.720 478.050 ;
        RECT 656.520 38.430 656.780 38.750 ;
        RECT 2851.640 38.430 2851.900 38.750 ;
        RECT 2851.700 2.400 2851.840 38.430 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
      LAYER via2 ;
        RECT 658.120 499.150 658.400 499.430 ;
        RECT 657.430 497.280 657.710 497.560 ;
      LAYER met3 ;
        RECT 658.095 499.125 658.425 499.455 ;
        RECT 657.405 497.570 657.735 497.585 ;
        RECT 658.110 497.570 658.410 499.125 ;
        RECT 657.405 497.270 658.410 497.570 ;
        RECT 657.405 497.255 657.735 497.270 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 659.480 499.500 659.800 499.760 ;
        RECT 659.570 498.400 659.710 499.500 ;
        RECT 659.250 498.200 659.710 498.400 ;
        RECT 659.250 498.140 659.570 498.200 ;
        RECT 657.410 473.520 657.730 473.580 ;
        RECT 659.250 473.520 659.570 473.580 ;
        RECT 657.410 473.380 659.570 473.520 ;
        RECT 657.410 473.320 657.730 473.380 ;
        RECT 659.250 473.320 659.570 473.380 ;
        RECT 657.410 38.320 657.730 38.380 ;
        RECT 2869.550 38.320 2869.870 38.380 ;
        RECT 657.410 38.180 2869.870 38.320 ;
        RECT 657.410 38.120 657.730 38.180 ;
        RECT 2869.550 38.120 2869.870 38.180 ;
      LAYER via ;
        RECT 659.510 499.500 659.770 499.760 ;
        RECT 659.280 498.140 659.540 498.400 ;
        RECT 657.440 473.320 657.700 473.580 ;
        RECT 659.280 473.320 659.540 473.580 ;
        RECT 657.440 38.120 657.700 38.380 ;
        RECT 2869.580 38.120 2869.840 38.380 ;
      LAYER met2 ;
        RECT 659.530 500.000 659.810 504.000 ;
        RECT 659.570 499.790 659.710 500.000 ;
        RECT 659.510 499.470 659.770 499.790 ;
        RECT 659.280 498.110 659.540 498.430 ;
        RECT 659.340 473.610 659.480 498.110 ;
        RECT 657.440 473.290 657.700 473.610 ;
        RECT 659.280 473.290 659.540 473.610 ;
        RECT 657.500 38.410 657.640 473.290 ;
        RECT 657.440 38.090 657.700 38.410 ;
        RECT 2869.580 38.090 2869.840 38.410 ;
        RECT 2869.640 2.400 2869.780 38.090 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 659.110 499.900 661.090 500.040 ;
        RECT 659.110 498.740 659.250 499.900 ;
        RECT 660.950 499.420 661.090 499.900 ;
        RECT 660.860 499.160 661.180 499.420 ;
        RECT 658.790 498.540 659.250 498.740 ;
        RECT 658.790 498.480 659.110 498.540 ;
      LAYER via ;
        RECT 660.890 499.160 661.150 499.420 ;
        RECT 658.820 498.480 659.080 498.740 ;
      LAYER met2 ;
        RECT 660.910 500.000 661.190 504.000 ;
        RECT 660.950 499.450 661.090 500.000 ;
        RECT 660.890 499.130 661.150 499.450 ;
        RECT 658.820 498.450 659.080 498.770 ;
        RECT 658.880 490.805 659.020 498.450 ;
        RECT 658.810 490.435 659.090 490.805 ;
        RECT 2884.290 120.515 2884.570 120.885 ;
        RECT 2884.360 82.870 2884.500 120.515 ;
        RECT 2884.360 82.730 2884.960 82.870 ;
        RECT 2884.820 1.770 2884.960 82.730 ;
        RECT 2886.910 1.770 2887.470 2.400 ;
        RECT 2884.820 1.630 2887.470 1.770 ;
        RECT 2886.910 -4.800 2887.470 1.630 ;
      LAYER via2 ;
        RECT 658.810 490.480 659.090 490.760 ;
        RECT 2884.290 120.560 2884.570 120.840 ;
      LAYER met3 ;
        RECT 658.070 490.770 658.450 490.780 ;
        RECT 658.785 490.770 659.115 490.785 ;
        RECT 658.070 490.470 659.115 490.770 ;
        RECT 658.070 490.460 658.450 490.470 ;
        RECT 658.785 490.455 659.115 490.470 ;
        RECT 658.070 120.850 658.450 120.860 ;
        RECT 2884.265 120.850 2884.595 120.865 ;
        RECT 658.070 120.550 2884.595 120.850 ;
        RECT 658.070 120.540 658.450 120.550 ;
        RECT 2884.265 120.535 2884.595 120.550 ;
      LAYER via3 ;
        RECT 658.100 490.460 658.420 490.780 ;
        RECT 658.100 120.540 658.420 120.860 ;
      LAYER met4 ;
        RECT 658.095 490.455 658.425 490.785 ;
        RECT 658.110 120.865 658.410 490.455 ;
        RECT 658.095 120.535 658.425 120.865 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 501.930 498.000 502.250 498.060 ;
        RECT 501.930 497.860 502.620 498.000 ;
        RECT 501.930 497.800 502.250 497.860 ;
        RECT 501.010 496.980 501.330 497.040 ;
        RECT 502.480 496.980 502.620 497.860 ;
        RECT 501.010 496.840 502.620 496.980 ;
        RECT 501.010 496.780 501.330 496.840 ;
        RECT 841.870 19.620 842.190 19.680 ;
        RECT 847.850 19.620 848.170 19.680 ;
        RECT 841.870 19.480 848.170 19.620 ;
        RECT 841.870 19.420 842.190 19.480 ;
        RECT 847.850 19.420 848.170 19.480 ;
      LAYER via ;
        RECT 501.960 497.800 502.220 498.060 ;
        RECT 501.040 496.780 501.300 497.040 ;
        RECT 841.900 19.420 842.160 19.680 ;
        RECT 847.880 19.420 848.140 19.680 ;
      LAYER met2 ;
        RECT 502.210 500.000 502.490 504.000 ;
        RECT 502.250 498.680 502.390 500.000 ;
        RECT 502.020 498.540 502.390 498.680 ;
        RECT 502.020 498.090 502.160 498.540 ;
        RECT 501.960 497.770 502.220 498.090 ;
        RECT 501.040 496.750 501.300 497.070 ;
        RECT 501.100 491.485 501.240 496.750 ;
        RECT 501.030 491.115 501.310 491.485 ;
        RECT 841.890 135.475 842.170 135.845 ;
        RECT 841.960 19.710 842.100 135.475 ;
        RECT 841.900 19.390 842.160 19.710 ;
        RECT 847.880 19.390 848.140 19.710 ;
        RECT 847.940 2.400 848.080 19.390 ;
        RECT 847.730 -4.800 848.290 2.400 ;
      LAYER via2 ;
        RECT 501.030 491.160 501.310 491.440 ;
        RECT 841.890 135.520 842.170 135.800 ;
      LAYER met3 ;
        RECT 501.005 491.460 501.335 491.465 ;
        RECT 500.750 491.450 501.335 491.460 ;
        RECT 500.550 491.150 501.335 491.450 ;
        RECT 500.750 491.140 501.335 491.150 ;
        RECT 501.005 491.135 501.335 491.140 ;
        RECT 500.750 135.810 501.130 135.820 ;
        RECT 841.865 135.810 842.195 135.825 ;
        RECT 500.750 135.510 842.195 135.810 ;
        RECT 500.750 135.500 501.130 135.510 ;
        RECT 841.865 135.495 842.195 135.510 ;
      LAYER via3 ;
        RECT 500.780 491.140 501.100 491.460 ;
        RECT 500.780 135.500 501.100 135.820 ;
      LAYER met4 ;
        RECT 500.775 491.135 501.105 491.465 ;
        RECT 500.790 135.825 501.090 491.135 ;
        RECT 500.775 135.495 501.105 135.825 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 503.310 490.520 503.630 490.580 ;
        RECT 504.230 490.520 504.550 490.580 ;
        RECT 503.310 490.380 504.550 490.520 ;
        RECT 503.310 490.320 503.630 490.380 ;
        RECT 504.230 490.320 504.550 490.380 ;
        RECT 504.230 473.520 504.550 473.580 ;
        RECT 505.150 473.520 505.470 473.580 ;
        RECT 504.230 473.380 505.470 473.520 ;
        RECT 504.230 473.320 504.550 473.380 ;
        RECT 505.150 473.320 505.470 473.380 ;
        RECT 505.150 122.640 505.470 122.700 ;
        RECT 862.570 122.640 862.890 122.700 ;
        RECT 505.150 122.500 862.890 122.640 ;
        RECT 505.150 122.440 505.470 122.500 ;
        RECT 862.570 122.440 862.890 122.500 ;
      LAYER via ;
        RECT 503.340 490.320 503.600 490.580 ;
        RECT 504.260 490.320 504.520 490.580 ;
        RECT 504.260 473.320 504.520 473.580 ;
        RECT 505.180 473.320 505.440 473.580 ;
        RECT 505.180 122.440 505.440 122.700 ;
        RECT 862.600 122.440 862.860 122.700 ;
      LAYER met2 ;
        RECT 503.590 500.000 503.870 504.000 ;
        RECT 503.630 498.340 503.770 500.000 ;
        RECT 503.400 498.200 503.770 498.340 ;
        RECT 503.400 490.610 503.540 498.200 ;
        RECT 503.340 490.290 503.600 490.610 ;
        RECT 504.260 490.290 504.520 490.610 ;
        RECT 504.320 473.610 504.460 490.290 ;
        RECT 504.260 473.290 504.520 473.610 ;
        RECT 505.180 473.290 505.440 473.610 ;
        RECT 505.240 122.730 505.380 473.290 ;
        RECT 505.180 122.410 505.440 122.730 ;
        RECT 862.600 122.410 862.860 122.730 ;
        RECT 862.660 82.870 862.800 122.410 ;
        RECT 862.660 82.730 863.720 82.870 ;
        RECT 863.580 1.770 863.720 82.730 ;
        RECT 865.670 1.770 866.230 2.400 ;
        RECT 863.580 1.630 866.230 1.770 ;
        RECT 865.670 -4.800 866.230 1.630 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.690 471.820 505.010 471.880 ;
        RECT 506.070 471.820 506.390 471.880 ;
        RECT 504.690 471.680 506.390 471.820 ;
        RECT 504.690 471.620 505.010 471.680 ;
        RECT 506.070 471.620 506.390 471.680 ;
        RECT 506.070 137.940 506.390 138.000 ;
        RECT 883.730 137.940 884.050 138.000 ;
        RECT 506.070 137.800 884.050 137.940 ;
        RECT 506.070 137.740 506.390 137.800 ;
        RECT 883.730 137.740 884.050 137.800 ;
      LAYER via ;
        RECT 504.720 471.620 504.980 471.880 ;
        RECT 506.100 471.620 506.360 471.880 ;
        RECT 506.100 137.740 506.360 138.000 ;
        RECT 883.760 137.740 884.020 138.000 ;
      LAYER met2 ;
        RECT 504.970 500.000 505.250 504.000 ;
        RECT 505.010 499.020 505.150 500.000 ;
        RECT 505.010 498.880 505.380 499.020 ;
        RECT 505.240 477.770 505.380 498.880 ;
        RECT 504.780 477.630 505.380 477.770 ;
        RECT 504.780 471.910 504.920 477.630 ;
        RECT 504.720 471.590 504.980 471.910 ;
        RECT 506.100 471.590 506.360 471.910 ;
        RECT 506.160 138.030 506.300 471.590 ;
        RECT 506.100 137.710 506.360 138.030 ;
        RECT 883.760 137.710 884.020 138.030 ;
        RECT 883.820 34.570 883.960 137.710 ;
        RECT 883.360 34.430 883.960 34.570 ;
        RECT 883.360 2.400 883.500 34.430 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 506.300 499.160 506.620 499.420 ;
        RECT 505.610 498.000 505.930 498.060 ;
        RECT 506.390 498.000 506.530 499.160 ;
        RECT 505.610 497.860 506.530 498.000 ;
        RECT 505.610 497.800 505.930 497.860 ;
        RECT 505.610 137.600 505.930 137.660 ;
        RECT 897.070 137.600 897.390 137.660 ;
        RECT 505.610 137.460 897.390 137.600 ;
        RECT 505.610 137.400 505.930 137.460 ;
        RECT 897.070 137.400 897.390 137.460 ;
      LAYER via ;
        RECT 506.330 499.160 506.590 499.420 ;
        RECT 505.640 497.800 505.900 498.060 ;
        RECT 505.640 137.400 505.900 137.660 ;
        RECT 897.100 137.400 897.360 137.660 ;
      LAYER met2 ;
        RECT 506.350 500.000 506.630 504.000 ;
        RECT 506.390 499.450 506.530 500.000 ;
        RECT 506.330 499.130 506.590 499.450 ;
        RECT 505.640 497.770 505.900 498.090 ;
        RECT 505.700 137.690 505.840 497.770 ;
        RECT 505.640 137.370 505.900 137.690 ;
        RECT 897.100 137.370 897.360 137.690 ;
        RECT 897.160 82.870 897.300 137.370 ;
        RECT 897.160 82.730 901.440 82.870 ;
        RECT 901.300 2.400 901.440 82.730 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 507.680 499.160 508.000 499.420 ;
        RECT 507.770 497.720 507.910 499.160 ;
        RECT 507.450 497.520 507.910 497.720 ;
        RECT 507.450 497.460 507.770 497.520 ;
        RECT 504.230 472.840 504.550 472.900 ;
        RECT 507.450 472.840 507.770 472.900 ;
        RECT 504.230 472.700 507.770 472.840 ;
        RECT 504.230 472.640 504.550 472.700 ;
        RECT 507.450 472.640 507.770 472.700 ;
        RECT 504.230 41.040 504.550 41.100 ;
        RECT 918.690 41.040 919.010 41.100 ;
        RECT 504.230 40.900 919.010 41.040 ;
        RECT 504.230 40.840 504.550 40.900 ;
        RECT 918.690 40.840 919.010 40.900 ;
      LAYER via ;
        RECT 507.710 499.160 507.970 499.420 ;
        RECT 507.480 497.460 507.740 497.720 ;
        RECT 504.260 472.640 504.520 472.900 ;
        RECT 507.480 472.640 507.740 472.900 ;
        RECT 504.260 40.840 504.520 41.100 ;
        RECT 918.720 40.840 918.980 41.100 ;
      LAYER met2 ;
        RECT 507.730 500.000 508.010 504.000 ;
        RECT 507.770 499.450 507.910 500.000 ;
        RECT 507.710 499.130 507.970 499.450 ;
        RECT 507.480 497.430 507.740 497.750 ;
        RECT 507.540 472.930 507.680 497.430 ;
        RECT 504.260 472.610 504.520 472.930 ;
        RECT 507.480 472.610 507.740 472.930 ;
        RECT 504.320 41.130 504.460 472.610 ;
        RECT 504.260 40.810 504.520 41.130 ;
        RECT 918.720 40.810 918.980 41.130 ;
        RECT 918.780 2.400 918.920 40.810 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 509.060 499.500 509.380 499.760 ;
        RECT 503.770 497.320 504.090 497.380 ;
        RECT 509.150 497.320 509.290 499.500 ;
        RECT 503.770 497.180 509.290 497.320 ;
        RECT 503.770 497.120 504.090 497.180 ;
        RECT 503.770 40.700 504.090 40.760 ;
        RECT 936.630 40.700 936.950 40.760 ;
        RECT 503.770 40.560 936.950 40.700 ;
        RECT 503.770 40.500 504.090 40.560 ;
        RECT 936.630 40.500 936.950 40.560 ;
      LAYER via ;
        RECT 509.090 499.500 509.350 499.760 ;
        RECT 503.800 497.120 504.060 497.380 ;
        RECT 503.800 40.500 504.060 40.760 ;
        RECT 936.660 40.500 936.920 40.760 ;
      LAYER met2 ;
        RECT 509.110 500.000 509.390 504.000 ;
        RECT 509.150 499.790 509.290 500.000 ;
        RECT 509.090 499.470 509.350 499.790 ;
        RECT 503.800 497.090 504.060 497.410 ;
        RECT 503.860 40.790 504.000 497.090 ;
        RECT 503.800 40.470 504.060 40.790 ;
        RECT 936.660 40.470 936.920 40.790 ;
        RECT 936.720 2.400 936.860 40.470 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.440 499.160 510.760 499.420 ;
        RECT 510.530 497.720 510.670 499.160 ;
        RECT 510.530 497.520 510.990 497.720 ;
        RECT 510.670 497.460 510.990 497.520 ;
        RECT 510.670 40.360 510.990 40.420 ;
        RECT 954.110 40.360 954.430 40.420 ;
        RECT 510.670 40.220 954.430 40.360 ;
        RECT 510.670 40.160 510.990 40.220 ;
        RECT 954.110 40.160 954.430 40.220 ;
      LAYER via ;
        RECT 510.470 499.160 510.730 499.420 ;
        RECT 510.700 497.460 510.960 497.720 ;
        RECT 510.700 40.160 510.960 40.420 ;
        RECT 954.140 40.160 954.400 40.420 ;
      LAYER met2 ;
        RECT 510.490 500.000 510.770 504.000 ;
        RECT 510.530 499.450 510.670 500.000 ;
        RECT 510.470 499.130 510.730 499.450 ;
        RECT 510.700 497.430 510.960 497.750 ;
        RECT 510.760 40.450 510.900 497.430 ;
        RECT 510.700 40.130 510.960 40.450 ;
        RECT 954.140 40.130 954.400 40.450 ;
        RECT 954.200 2.400 954.340 40.130 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.820 499.160 512.140 499.420 ;
        RECT 511.910 497.660 512.050 499.160 ;
        RECT 512.510 497.660 512.830 497.720 ;
        RECT 511.910 497.520 512.830 497.660 ;
        RECT 512.510 497.460 512.830 497.520 ;
        RECT 512.510 122.300 512.830 122.360 ;
        RECT 966.070 122.300 966.390 122.360 ;
        RECT 512.510 122.160 966.390 122.300 ;
        RECT 512.510 122.100 512.830 122.160 ;
        RECT 966.070 122.100 966.390 122.160 ;
        RECT 966.070 19.620 966.390 19.680 ;
        RECT 972.050 19.620 972.370 19.680 ;
        RECT 966.070 19.480 972.370 19.620 ;
        RECT 966.070 19.420 966.390 19.480 ;
        RECT 972.050 19.420 972.370 19.480 ;
      LAYER via ;
        RECT 511.850 499.160 512.110 499.420 ;
        RECT 512.540 497.460 512.800 497.720 ;
        RECT 512.540 122.100 512.800 122.360 ;
        RECT 966.100 122.100 966.360 122.360 ;
        RECT 966.100 19.420 966.360 19.680 ;
        RECT 972.080 19.420 972.340 19.680 ;
      LAYER met2 ;
        RECT 511.870 500.000 512.150 504.000 ;
        RECT 511.910 499.450 512.050 500.000 ;
        RECT 511.850 499.130 512.110 499.450 ;
        RECT 512.540 497.430 512.800 497.750 ;
        RECT 512.600 122.390 512.740 497.430 ;
        RECT 512.540 122.070 512.800 122.390 ;
        RECT 966.100 122.070 966.360 122.390 ;
        RECT 966.160 19.710 966.300 122.070 ;
        RECT 966.100 19.390 966.360 19.710 ;
        RECT 972.080 19.390 972.340 19.710 ;
        RECT 972.140 2.400 972.280 19.390 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 484.450 472.840 484.770 472.900 ;
        RECT 486.750 472.840 487.070 472.900 ;
        RECT 484.450 472.700 487.070 472.840 ;
        RECT 484.450 472.640 484.770 472.700 ;
        RECT 486.750 472.640 487.070 472.700 ;
        RECT 541.950 18.260 542.270 18.320 ;
        RECT 652.810 18.260 653.130 18.320 ;
        RECT 541.950 18.120 653.130 18.260 ;
        RECT 541.950 18.060 542.270 18.120 ;
        RECT 652.810 18.060 653.130 18.120 ;
        RECT 484.450 16.220 484.770 16.280 ;
        RECT 541.950 16.220 542.270 16.280 ;
        RECT 484.450 16.080 542.270 16.220 ;
        RECT 484.450 16.020 484.770 16.080 ;
        RECT 541.950 16.020 542.270 16.080 ;
      LAYER via ;
        RECT 484.480 472.640 484.740 472.900 ;
        RECT 486.780 472.640 487.040 472.900 ;
        RECT 541.980 18.060 542.240 18.320 ;
        RECT 652.840 18.060 653.100 18.320 ;
        RECT 484.480 16.020 484.740 16.280 ;
        RECT 541.980 16.020 542.240 16.280 ;
      LAYER met2 ;
        RECT 487.030 500.000 487.310 504.000 ;
        RECT 487.070 498.340 487.210 500.000 ;
        RECT 486.840 498.200 487.210 498.340 ;
        RECT 486.840 472.930 486.980 498.200 ;
        RECT 484.480 472.610 484.740 472.930 ;
        RECT 486.780 472.610 487.040 472.930 ;
        RECT 484.540 16.310 484.680 472.610 ;
        RECT 541.980 18.030 542.240 18.350 ;
        RECT 652.840 18.030 653.100 18.350 ;
        RECT 542.040 16.310 542.180 18.030 ;
        RECT 484.480 15.990 484.740 16.310 ;
        RECT 541.980 15.990 542.240 16.310 ;
        RECT 652.900 2.400 653.040 18.030 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 512.970 137.260 513.290 137.320 ;
        RECT 986.770 137.260 987.090 137.320 ;
        RECT 512.970 137.120 987.090 137.260 ;
        RECT 512.970 137.060 513.290 137.120 ;
        RECT 986.770 137.060 987.090 137.120 ;
      LAYER via ;
        RECT 513.000 137.060 513.260 137.320 ;
        RECT 986.800 137.060 987.060 137.320 ;
      LAYER met2 ;
        RECT 513.250 500.000 513.530 504.000 ;
        RECT 513.290 498.340 513.430 500.000 ;
        RECT 513.060 498.200 513.430 498.340 ;
        RECT 513.060 137.350 513.200 498.200 ;
        RECT 513.000 137.030 513.260 137.350 ;
        RECT 986.800 137.030 987.060 137.350 ;
        RECT 986.860 82.870 987.000 137.030 ;
        RECT 986.860 82.730 989.760 82.870 ;
        RECT 989.620 2.400 989.760 82.730 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.630 500.000 514.910 504.000 ;
        RECT 514.670 498.680 514.810 500.000 ;
        RECT 514.440 498.540 514.810 498.680 ;
        RECT 514.440 483.325 514.580 498.540 ;
        RECT 514.370 482.955 514.650 483.325 ;
        RECT 1007.950 143.635 1008.230 144.005 ;
        RECT 1008.020 34.570 1008.160 143.635 ;
        RECT 1007.560 34.430 1008.160 34.570 ;
        RECT 1007.560 2.400 1007.700 34.430 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
      LAYER via2 ;
        RECT 514.370 483.000 514.650 483.280 ;
        RECT 1007.950 143.680 1008.230 143.960 ;
      LAYER met3 ;
        RECT 514.345 483.300 514.675 483.305 ;
        RECT 514.345 483.290 514.930 483.300 ;
        RECT 514.120 482.990 514.930 483.290 ;
        RECT 514.345 482.980 514.930 482.990 ;
        RECT 514.345 482.975 514.675 482.980 ;
        RECT 514.550 143.970 514.930 143.980 ;
        RECT 1007.925 143.970 1008.255 143.985 ;
        RECT 514.550 143.670 1008.255 143.970 ;
        RECT 514.550 143.660 514.930 143.670 ;
        RECT 1007.925 143.655 1008.255 143.670 ;
      LAYER via3 ;
        RECT 514.580 482.980 514.900 483.300 ;
        RECT 514.580 143.660 514.900 143.980 ;
      LAYER met4 ;
        RECT 514.575 482.975 514.905 483.305 ;
        RECT 514.590 143.985 514.890 482.975 ;
        RECT 514.575 143.655 514.905 143.985 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 516.190 490.860 516.510 490.920 ;
        RECT 524.010 490.860 524.330 490.920 ;
        RECT 516.190 490.720 524.330 490.860 ;
        RECT 516.190 490.660 516.510 490.720 ;
        RECT 524.010 490.660 524.330 490.720 ;
        RECT 524.010 485.760 524.330 485.820 ;
        RECT 543.790 485.760 544.110 485.820 ;
        RECT 524.010 485.620 544.110 485.760 ;
        RECT 524.010 485.560 524.330 485.620 ;
        RECT 543.790 485.560 544.110 485.620 ;
        RECT 542.870 143.720 543.190 143.780 ;
        RECT 1021.270 143.720 1021.590 143.780 ;
        RECT 542.870 143.580 1021.590 143.720 ;
        RECT 542.870 143.520 543.190 143.580 ;
        RECT 1021.270 143.520 1021.590 143.580 ;
      LAYER via ;
        RECT 516.220 490.660 516.480 490.920 ;
        RECT 524.040 490.660 524.300 490.920 ;
        RECT 524.040 485.560 524.300 485.820 ;
        RECT 543.820 485.560 544.080 485.820 ;
        RECT 542.900 143.520 543.160 143.780 ;
        RECT 1021.300 143.520 1021.560 143.780 ;
      LAYER met2 ;
        RECT 516.010 500.000 516.290 504.000 ;
        RECT 516.050 498.340 516.190 500.000 ;
        RECT 516.050 498.200 516.420 498.340 ;
        RECT 516.280 490.950 516.420 498.200 ;
        RECT 516.220 490.630 516.480 490.950 ;
        RECT 524.040 490.630 524.300 490.950 ;
        RECT 524.100 485.850 524.240 490.630 ;
        RECT 524.040 485.530 524.300 485.850 ;
        RECT 543.820 485.530 544.080 485.850 ;
        RECT 543.880 448.570 544.020 485.530 ;
        RECT 542.960 448.430 544.020 448.570 ;
        RECT 542.960 143.810 543.100 448.430 ;
        RECT 542.900 143.490 543.160 143.810 ;
        RECT 1021.300 143.490 1021.560 143.810 ;
        RECT 1021.360 82.870 1021.500 143.490 ;
        RECT 1021.360 82.730 1025.640 82.870 ;
        RECT 1025.500 2.400 1025.640 82.730 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.340 499.500 517.660 499.760 ;
        RECT 517.430 499.080 517.570 499.500 ;
        RECT 517.110 498.880 517.570 499.080 ;
        RECT 517.110 498.820 517.430 498.880 ;
        RECT 517.110 490.180 517.430 490.240 ;
        RECT 518.490 490.180 518.810 490.240 ;
        RECT 517.110 490.040 518.810 490.180 ;
        RECT 517.110 489.980 517.430 490.040 ;
        RECT 518.490 489.980 518.810 490.040 ;
        RECT 518.950 47.160 519.270 47.220 ;
        RECT 1042.890 47.160 1043.210 47.220 ;
        RECT 518.950 47.020 1043.210 47.160 ;
        RECT 518.950 46.960 519.270 47.020 ;
        RECT 1042.890 46.960 1043.210 47.020 ;
      LAYER via ;
        RECT 517.370 499.500 517.630 499.760 ;
        RECT 517.140 498.820 517.400 499.080 ;
        RECT 517.140 489.980 517.400 490.240 ;
        RECT 518.520 489.980 518.780 490.240 ;
        RECT 518.980 46.960 519.240 47.220 ;
        RECT 1042.920 46.960 1043.180 47.220 ;
      LAYER met2 ;
        RECT 517.390 500.000 517.670 504.000 ;
        RECT 517.430 499.790 517.570 500.000 ;
        RECT 517.370 499.470 517.630 499.790 ;
        RECT 517.140 498.790 517.400 499.110 ;
        RECT 517.200 490.270 517.340 498.790 ;
        RECT 517.140 489.950 517.400 490.270 ;
        RECT 518.520 489.950 518.780 490.270 ;
        RECT 518.580 481.170 518.720 489.950 ;
        RECT 518.580 481.030 519.180 481.170 ;
        RECT 519.040 47.250 519.180 481.030 ;
        RECT 518.980 46.930 519.240 47.250 ;
        RECT 1042.920 46.930 1043.180 47.250 ;
        RECT 1042.980 2.400 1043.120 46.930 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.030 46.820 518.350 46.880 ;
        RECT 1060.830 46.820 1061.150 46.880 ;
        RECT 518.030 46.680 1061.150 46.820 ;
        RECT 518.030 46.620 518.350 46.680 ;
        RECT 1060.830 46.620 1061.150 46.680 ;
      LAYER via ;
        RECT 518.060 46.620 518.320 46.880 ;
        RECT 1060.860 46.620 1061.120 46.880 ;
      LAYER met2 ;
        RECT 518.770 500.000 519.050 504.000 ;
        RECT 518.810 498.680 518.950 500.000 ;
        RECT 518.580 498.540 518.950 498.680 ;
        RECT 518.580 492.050 518.720 498.540 ;
        RECT 518.120 491.910 518.720 492.050 ;
        RECT 518.120 46.910 518.260 491.910 ;
        RECT 518.060 46.590 518.320 46.910 ;
        RECT 1060.860 46.590 1061.120 46.910 ;
        RECT 1060.920 2.400 1061.060 46.590 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.810 499.900 520.330 500.040 ;
        RECT 518.810 497.040 518.950 499.900 ;
        RECT 520.190 499.760 520.330 499.900 ;
        RECT 520.100 499.500 520.420 499.760 ;
        RECT 518.810 496.840 519.270 497.040 ;
        RECT 518.950 496.780 519.270 496.840 ;
        RECT 518.950 481.480 519.270 481.740 ;
        RECT 518.490 480.660 518.810 480.720 ;
        RECT 519.040 480.660 519.180 481.480 ;
        RECT 518.490 480.520 519.180 480.660 ;
        RECT 518.490 480.460 518.810 480.520 ;
        RECT 518.490 46.480 518.810 46.540 ;
        RECT 1078.310 46.480 1078.630 46.540 ;
        RECT 518.490 46.340 1078.630 46.480 ;
        RECT 518.490 46.280 518.810 46.340 ;
        RECT 1078.310 46.280 1078.630 46.340 ;
      LAYER via ;
        RECT 520.130 499.500 520.390 499.760 ;
        RECT 518.980 496.780 519.240 497.040 ;
        RECT 518.980 481.480 519.240 481.740 ;
        RECT 518.520 480.460 518.780 480.720 ;
        RECT 518.520 46.280 518.780 46.540 ;
        RECT 1078.340 46.280 1078.600 46.540 ;
      LAYER met2 ;
        RECT 520.150 500.000 520.430 504.000 ;
        RECT 520.190 499.790 520.330 500.000 ;
        RECT 520.130 499.470 520.390 499.790 ;
        RECT 518.980 496.750 519.240 497.070 ;
        RECT 519.040 481.770 519.180 496.750 ;
        RECT 518.980 481.450 519.240 481.770 ;
        RECT 518.520 480.430 518.780 480.750 ;
        RECT 518.580 46.570 518.720 480.430 ;
        RECT 518.520 46.250 518.780 46.570 ;
        RECT 1078.340 46.250 1078.600 46.570 ;
        RECT 1078.400 2.400 1078.540 46.250 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 521.250 483.720 521.570 483.780 ;
        RECT 521.250 483.580 531.370 483.720 ;
        RECT 521.250 483.520 521.570 483.580 ;
        RECT 531.230 483.380 531.370 483.580 ;
        RECT 557.130 483.380 557.450 483.440 ;
        RECT 531.230 483.240 557.450 483.380 ;
        RECT 557.130 483.180 557.450 483.240 ;
        RECT 557.130 143.380 557.450 143.440 ;
        RECT 1090.270 143.380 1090.590 143.440 ;
        RECT 557.130 143.240 1090.590 143.380 ;
        RECT 557.130 143.180 557.450 143.240 ;
        RECT 1090.270 143.180 1090.590 143.240 ;
        RECT 1090.270 58.380 1090.590 58.440 ;
        RECT 1096.250 58.380 1096.570 58.440 ;
        RECT 1090.270 58.240 1096.570 58.380 ;
        RECT 1090.270 58.180 1090.590 58.240 ;
        RECT 1096.250 58.180 1096.570 58.240 ;
      LAYER via ;
        RECT 521.280 483.520 521.540 483.780 ;
        RECT 557.160 483.180 557.420 483.440 ;
        RECT 557.160 143.180 557.420 143.440 ;
        RECT 1090.300 143.180 1090.560 143.440 ;
        RECT 1090.300 58.180 1090.560 58.440 ;
        RECT 1096.280 58.180 1096.540 58.440 ;
      LAYER met2 ;
        RECT 521.530 500.000 521.810 504.000 ;
        RECT 521.570 498.340 521.710 500.000 ;
        RECT 521.340 498.200 521.710 498.340 ;
        RECT 521.340 483.810 521.480 498.200 ;
        RECT 521.280 483.490 521.540 483.810 ;
        RECT 557.160 483.150 557.420 483.470 ;
        RECT 557.220 143.470 557.360 483.150 ;
        RECT 557.160 143.150 557.420 143.470 ;
        RECT 1090.300 143.150 1090.560 143.470 ;
        RECT 1090.360 58.470 1090.500 143.150 ;
        RECT 1090.300 58.150 1090.560 58.470 ;
        RECT 1096.280 58.150 1096.540 58.470 ;
        RECT 1096.340 2.400 1096.480 58.150 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.910 500.000 523.190 504.000 ;
        RECT 522.950 499.135 523.090 500.000 ;
        RECT 522.880 498.765 523.160 499.135 ;
        RECT 1113.750 52.515 1114.030 52.885 ;
        RECT 1113.820 2.400 1113.960 52.515 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
      LAYER via2 ;
        RECT 522.880 498.810 523.160 499.090 ;
        RECT 1113.750 52.560 1114.030 52.840 ;
      LAYER met3 ;
        RECT 522.855 498.930 523.185 499.115 ;
        RECT 523.750 498.930 524.130 498.940 ;
        RECT 522.855 498.785 524.130 498.930 ;
        RECT 522.870 498.630 524.130 498.785 ;
        RECT 523.750 498.620 524.130 498.630 ;
        RECT 523.750 52.850 524.130 52.860 ;
        RECT 1113.725 52.850 1114.055 52.865 ;
        RECT 523.750 52.550 1114.055 52.850 ;
        RECT 523.750 52.540 524.130 52.550 ;
        RECT 1113.725 52.535 1114.055 52.550 ;
      LAYER via3 ;
        RECT 523.780 498.620 524.100 498.940 ;
        RECT 523.780 52.540 524.100 52.860 ;
      LAYER met4 ;
        RECT 523.775 498.615 524.105 498.945 ;
        RECT 523.790 52.865 524.090 498.615 ;
        RECT 523.775 52.535 524.105 52.865 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.240 499.500 524.560 499.760 ;
        RECT 524.330 498.740 524.470 499.500 ;
        RECT 524.010 498.540 524.470 498.740 ;
        RECT 524.010 498.480 524.330 498.540 ;
        RECT 524.930 46.140 525.250 46.200 ;
        RECT 1132.130 46.140 1132.450 46.200 ;
        RECT 524.930 46.000 1132.450 46.140 ;
        RECT 524.930 45.940 525.250 46.000 ;
        RECT 1132.130 45.940 1132.450 46.000 ;
      LAYER via ;
        RECT 524.270 499.500 524.530 499.760 ;
        RECT 524.040 498.480 524.300 498.740 ;
        RECT 524.960 45.940 525.220 46.200 ;
        RECT 1132.160 45.940 1132.420 46.200 ;
      LAYER met2 ;
        RECT 524.290 500.000 524.570 504.000 ;
        RECT 524.330 499.790 524.470 500.000 ;
        RECT 524.270 499.470 524.530 499.790 ;
        RECT 524.040 498.450 524.300 498.770 ;
        RECT 524.100 491.540 524.240 498.450 ;
        RECT 524.100 491.400 525.160 491.540 ;
        RECT 525.020 46.230 525.160 491.400 ;
        RECT 524.960 45.910 525.220 46.230 ;
        RECT 1132.160 45.910 1132.420 46.230 ;
        RECT 1132.220 17.410 1132.360 45.910 ;
        RECT 1131.760 17.270 1132.360 17.410 ;
        RECT 1131.760 2.400 1131.900 17.270 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 525.620 499.500 525.940 499.760 ;
        RECT 525.710 498.400 525.850 499.500 ;
        RECT 525.390 498.200 525.850 498.400 ;
        RECT 525.390 498.140 525.710 498.200 ;
        RECT 525.390 53.280 525.710 53.340 ;
        RECT 1146.850 53.280 1147.170 53.340 ;
        RECT 525.390 53.140 1147.170 53.280 ;
        RECT 525.390 53.080 525.710 53.140 ;
        RECT 1146.850 53.080 1147.170 53.140 ;
      LAYER via ;
        RECT 525.650 499.500 525.910 499.760 ;
        RECT 525.420 498.140 525.680 498.400 ;
        RECT 525.420 53.080 525.680 53.340 ;
        RECT 1146.880 53.080 1147.140 53.340 ;
      LAYER met2 ;
        RECT 525.670 500.000 525.950 504.000 ;
        RECT 525.710 499.790 525.850 500.000 ;
        RECT 525.650 499.470 525.910 499.790 ;
        RECT 525.420 498.110 525.680 498.430 ;
        RECT 525.480 53.370 525.620 498.110 ;
        RECT 525.420 53.050 525.680 53.370 ;
        RECT 1146.880 53.050 1147.140 53.370 ;
        RECT 1146.940 1.770 1147.080 53.050 ;
        RECT 1149.030 1.770 1149.590 2.400 ;
        RECT 1146.940 1.630 1149.590 1.770 ;
        RECT 1149.030 -4.800 1149.590 1.630 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.410 500.000 488.690 504.000 ;
        RECT 488.450 499.645 488.590 500.000 ;
        RECT 488.380 499.275 488.660 499.645 ;
        RECT 670.770 27.355 671.050 27.725 ;
        RECT 670.840 2.400 670.980 27.355 ;
        RECT 670.630 -4.800 671.190 2.400 ;
      LAYER via2 ;
        RECT 488.380 499.320 488.660 499.600 ;
        RECT 670.770 27.400 671.050 27.680 ;
      LAYER met3 ;
        RECT 488.355 499.610 488.685 499.625 ;
        RECT 488.355 499.295 488.900 499.610 ;
        RECT 487.870 498.930 488.250 498.940 ;
        RECT 488.600 498.930 488.900 499.295 ;
        RECT 487.870 498.630 488.900 498.930 ;
        RECT 487.870 498.620 488.250 498.630 ;
        RECT 487.870 27.690 488.250 27.700 ;
        RECT 670.745 27.690 671.075 27.705 ;
        RECT 487.870 27.390 671.075 27.690 ;
        RECT 487.870 27.380 488.250 27.390 ;
        RECT 670.745 27.375 671.075 27.390 ;
      LAYER via3 ;
        RECT 487.900 498.620 488.220 498.940 ;
        RECT 487.900 27.380 488.220 27.700 ;
      LAYER met4 ;
        RECT 487.895 498.615 488.225 498.945 ;
        RECT 487.910 27.705 488.210 498.615 ;
        RECT 487.895 27.375 488.225 27.705 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.000 499.160 527.320 499.420 ;
        RECT 527.090 498.060 527.230 499.160 ;
        RECT 527.090 497.860 527.550 498.060 ;
        RECT 527.230 497.800 527.550 497.860 ;
        RECT 526.770 121.960 527.090 122.020 ;
        RECT 1166.170 121.960 1166.490 122.020 ;
        RECT 526.770 121.820 1166.490 121.960 ;
        RECT 526.770 121.760 527.090 121.820 ;
        RECT 1166.170 121.760 1166.490 121.820 ;
      LAYER via ;
        RECT 527.030 499.160 527.290 499.420 ;
        RECT 527.260 497.800 527.520 498.060 ;
        RECT 526.800 121.760 527.060 122.020 ;
        RECT 1166.200 121.760 1166.460 122.020 ;
      LAYER met2 ;
        RECT 527.050 500.000 527.330 504.000 ;
        RECT 527.090 499.450 527.230 500.000 ;
        RECT 527.030 499.130 527.290 499.450 ;
        RECT 527.260 497.770 527.520 498.090 ;
        RECT 527.320 488.650 527.460 497.770 ;
        RECT 526.860 488.510 527.460 488.650 ;
        RECT 526.860 122.050 527.000 488.510 ;
        RECT 526.800 121.730 527.060 122.050 ;
        RECT 1166.200 121.730 1166.460 122.050 ;
        RECT 1166.260 82.870 1166.400 121.730 ;
        RECT 1166.260 82.730 1167.320 82.870 ;
        RECT 1167.180 2.400 1167.320 82.730 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 528.380 498.820 528.700 499.080 ;
        RECT 528.470 498.680 528.610 498.820 ;
        RECT 528.470 498.540 528.840 498.680 ;
        RECT 527.690 498.000 528.010 498.060 ;
        RECT 528.700 498.000 528.840 498.540 ;
        RECT 527.690 497.860 528.840 498.000 ;
        RECT 527.690 497.800 528.010 497.860 ;
        RECT 525.850 473.520 526.170 473.580 ;
        RECT 527.690 473.520 528.010 473.580 ;
        RECT 525.850 473.380 528.010 473.520 ;
        RECT 525.850 473.320 526.170 473.380 ;
        RECT 527.690 473.320 528.010 473.380 ;
        RECT 525.850 52.940 526.170 53.000 ;
        RECT 1182.730 52.940 1183.050 53.000 ;
        RECT 525.850 52.800 1183.050 52.940 ;
        RECT 525.850 52.740 526.170 52.800 ;
        RECT 1182.730 52.740 1183.050 52.800 ;
      LAYER via ;
        RECT 528.410 498.820 528.670 499.080 ;
        RECT 527.720 497.800 527.980 498.060 ;
        RECT 525.880 473.320 526.140 473.580 ;
        RECT 527.720 473.320 527.980 473.580 ;
        RECT 525.880 52.740 526.140 53.000 ;
        RECT 1182.760 52.740 1183.020 53.000 ;
      LAYER met2 ;
        RECT 528.430 500.000 528.710 504.000 ;
        RECT 528.470 499.110 528.610 500.000 ;
        RECT 528.410 498.790 528.670 499.110 ;
        RECT 527.720 497.770 527.980 498.090 ;
        RECT 527.780 473.610 527.920 497.770 ;
        RECT 525.880 473.290 526.140 473.610 ;
        RECT 527.720 473.290 527.980 473.610 ;
        RECT 525.940 53.030 526.080 473.290 ;
        RECT 525.880 52.710 526.140 53.030 ;
        RECT 1182.760 52.710 1183.020 53.030 ;
        RECT 1182.820 1.770 1182.960 52.710 ;
        RECT 1184.910 1.770 1185.470 2.400 ;
        RECT 1182.820 1.630 1185.470 1.770 ;
        RECT 1184.910 -4.800 1185.470 1.630 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.810 500.000 530.090 504.000 ;
        RECT 529.850 499.645 529.990 500.000 ;
        RECT 529.780 499.275 530.060 499.645 ;
        RECT 1200.690 142.955 1200.970 143.325 ;
        RECT 1200.760 1.770 1200.900 142.955 ;
        RECT 1202.390 1.770 1202.950 2.400 ;
        RECT 1200.760 1.630 1202.950 1.770 ;
        RECT 1202.390 -4.800 1202.950 1.630 ;
      LAYER via2 ;
        RECT 529.780 499.320 530.060 499.600 ;
        RECT 1200.690 143.000 1200.970 143.280 ;
      LAYER met3 ;
        RECT 525.590 499.610 525.970 499.620 ;
        RECT 529.755 499.610 530.085 499.625 ;
        RECT 525.590 499.310 530.085 499.610 ;
        RECT 525.590 499.300 525.970 499.310 ;
        RECT 529.755 499.295 530.085 499.310 ;
        RECT 525.590 143.290 525.970 143.300 ;
        RECT 1200.665 143.290 1200.995 143.305 ;
        RECT 525.590 142.990 1200.995 143.290 ;
        RECT 525.590 142.980 525.970 142.990 ;
        RECT 1200.665 142.975 1200.995 142.990 ;
      LAYER via3 ;
        RECT 525.620 499.300 525.940 499.620 ;
        RECT 525.620 142.980 525.940 143.300 ;
      LAYER met4 ;
        RECT 525.615 499.295 525.945 499.625 ;
        RECT 525.630 143.305 525.930 499.295 ;
        RECT 525.615 142.975 525.945 143.305 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.370 477.600 531.690 477.660 ;
        RECT 534.130 477.600 534.450 477.660 ;
        RECT 531.370 477.460 534.450 477.600 ;
        RECT 531.370 477.400 531.690 477.460 ;
        RECT 534.130 477.400 534.450 477.460 ;
        RECT 534.130 143.040 534.450 143.100 ;
        RECT 1214.470 143.040 1214.790 143.100 ;
        RECT 534.130 142.900 1214.790 143.040 ;
        RECT 534.130 142.840 534.450 142.900 ;
        RECT 1214.470 142.840 1214.790 142.900 ;
        RECT 1214.470 58.380 1214.790 58.440 ;
        RECT 1220.450 58.380 1220.770 58.440 ;
        RECT 1214.470 58.240 1220.770 58.380 ;
        RECT 1214.470 58.180 1214.790 58.240 ;
        RECT 1220.450 58.180 1220.770 58.240 ;
      LAYER via ;
        RECT 531.400 477.400 531.660 477.660 ;
        RECT 534.160 477.400 534.420 477.660 ;
        RECT 534.160 142.840 534.420 143.100 ;
        RECT 1214.500 142.840 1214.760 143.100 ;
        RECT 1214.500 58.180 1214.760 58.440 ;
        RECT 1220.480 58.180 1220.740 58.440 ;
      LAYER met2 ;
        RECT 531.190 500.000 531.470 504.000 ;
        RECT 531.230 498.000 531.370 500.000 ;
        RECT 531.230 497.860 531.600 498.000 ;
        RECT 531.460 477.690 531.600 497.860 ;
        RECT 531.400 477.370 531.660 477.690 ;
        RECT 534.160 477.370 534.420 477.690 ;
        RECT 534.220 143.130 534.360 477.370 ;
        RECT 534.160 142.810 534.420 143.130 ;
        RECT 1214.500 142.810 1214.760 143.130 ;
        RECT 1214.560 58.470 1214.700 142.810 ;
        RECT 1214.500 58.150 1214.760 58.470 ;
        RECT 1220.480 58.150 1220.740 58.470 ;
        RECT 1220.540 2.400 1220.680 58.150 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 532.520 499.500 532.840 499.760 ;
        RECT 532.610 498.400 532.750 499.500 ;
        RECT 532.610 498.200 533.070 498.400 ;
        RECT 532.750 498.140 533.070 498.200 ;
        RECT 532.290 52.600 532.610 52.660 ;
        RECT 1237.930 52.600 1238.250 52.660 ;
        RECT 532.290 52.460 1238.250 52.600 ;
        RECT 532.290 52.400 532.610 52.460 ;
        RECT 1237.930 52.400 1238.250 52.460 ;
      LAYER via ;
        RECT 532.550 499.500 532.810 499.760 ;
        RECT 532.780 498.140 533.040 498.400 ;
        RECT 532.320 52.400 532.580 52.660 ;
        RECT 1237.960 52.400 1238.220 52.660 ;
      LAYER met2 ;
        RECT 532.570 500.000 532.850 504.000 ;
        RECT 532.610 499.790 532.750 500.000 ;
        RECT 532.550 499.470 532.810 499.790 ;
        RECT 532.780 498.110 533.040 498.430 ;
        RECT 532.840 488.140 532.980 498.110 ;
        RECT 532.380 488.000 532.980 488.140 ;
        RECT 532.380 52.690 532.520 488.000 ;
        RECT 532.320 52.370 532.580 52.690 ;
        RECT 1237.960 52.370 1238.220 52.690 ;
        RECT 1238.020 2.400 1238.160 52.370 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.830 52.260 532.150 52.320 ;
        RECT 1256.330 52.260 1256.650 52.320 ;
        RECT 531.830 52.120 1256.650 52.260 ;
        RECT 531.830 52.060 532.150 52.120 ;
        RECT 1256.330 52.060 1256.650 52.120 ;
      LAYER via ;
        RECT 531.860 52.060 532.120 52.320 ;
        RECT 1256.360 52.060 1256.620 52.320 ;
      LAYER met2 ;
        RECT 533.950 500.000 534.230 504.000 ;
        RECT 533.990 499.815 534.130 500.000 ;
        RECT 533.920 499.445 534.200 499.815 ;
        RECT 532.310 497.235 532.590 497.605 ;
        RECT 532.380 488.650 532.520 497.235 ;
        RECT 531.920 488.510 532.520 488.650 ;
        RECT 531.920 52.350 532.060 488.510 ;
        RECT 531.860 52.030 532.120 52.350 ;
        RECT 1256.360 52.030 1256.620 52.350 ;
        RECT 1256.420 17.410 1256.560 52.030 ;
        RECT 1255.960 17.270 1256.560 17.410 ;
        RECT 1255.960 2.400 1256.100 17.270 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
      LAYER via2 ;
        RECT 533.920 499.490 534.200 499.770 ;
        RECT 532.310 497.280 532.590 497.560 ;
      LAYER met3 ;
        RECT 533.895 499.465 534.225 499.795 ;
        RECT 532.285 497.570 532.615 497.585 ;
        RECT 533.910 497.570 534.210 499.465 ;
        RECT 532.285 497.270 534.210 497.570 ;
        RECT 532.285 497.255 532.615 497.270 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 535.280 499.500 535.600 499.760 ;
        RECT 535.370 498.400 535.510 499.500 ;
        RECT 535.370 498.200 535.830 498.400 ;
        RECT 535.510 498.140 535.830 498.200 ;
        RECT 532.750 487.460 533.070 487.520 ;
        RECT 535.510 487.460 535.830 487.520 ;
        RECT 532.750 487.320 535.830 487.460 ;
        RECT 532.750 487.260 533.070 487.320 ;
        RECT 535.510 487.260 535.830 487.320 ;
        RECT 532.750 60.080 533.070 60.140 ;
        RECT 1271.050 60.080 1271.370 60.140 ;
        RECT 532.750 59.940 1271.370 60.080 ;
        RECT 532.750 59.880 533.070 59.940 ;
        RECT 1271.050 59.880 1271.370 59.940 ;
      LAYER via ;
        RECT 535.310 499.500 535.570 499.760 ;
        RECT 535.540 498.140 535.800 498.400 ;
        RECT 532.780 487.260 533.040 487.520 ;
        RECT 535.540 487.260 535.800 487.520 ;
        RECT 532.780 59.880 533.040 60.140 ;
        RECT 1271.080 59.880 1271.340 60.140 ;
      LAYER met2 ;
        RECT 535.330 500.000 535.610 504.000 ;
        RECT 535.370 499.790 535.510 500.000 ;
        RECT 535.310 499.470 535.570 499.790 ;
        RECT 535.540 498.110 535.800 498.430 ;
        RECT 535.600 487.550 535.740 498.110 ;
        RECT 532.780 487.230 533.040 487.550 ;
        RECT 535.540 487.230 535.800 487.550 ;
        RECT 532.840 60.170 532.980 487.230 ;
        RECT 532.780 59.850 533.040 60.170 ;
        RECT 1271.080 59.850 1271.340 60.170 ;
        RECT 1271.140 1.770 1271.280 59.850 ;
        RECT 1273.230 1.770 1273.790 2.400 ;
        RECT 1271.140 1.630 1273.790 1.770 ;
        RECT 1273.230 -4.800 1273.790 1.630 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 536.660 500.860 536.980 501.120 ;
        RECT 536.750 499.020 536.890 500.860 ;
        RECT 536.750 498.880 537.580 499.020 ;
        RECT 537.440 498.400 537.580 498.880 ;
        RECT 537.350 498.140 537.670 498.400 ;
      LAYER via ;
        RECT 536.690 500.860 536.950 501.120 ;
        RECT 537.380 498.140 537.640 498.400 ;
      LAYER met2 ;
        RECT 536.710 501.150 536.990 504.000 ;
        RECT 536.690 500.830 536.990 501.150 ;
        RECT 536.710 500.000 536.990 500.830 ;
        RECT 537.380 498.110 537.640 498.430 ;
        RECT 537.440 492.165 537.580 498.110 ;
        RECT 537.370 491.795 537.650 492.165 ;
        RECT 1291.310 59.315 1291.590 59.685 ;
        RECT 1291.380 2.400 1291.520 59.315 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
      LAYER via2 ;
        RECT 537.370 491.840 537.650 492.120 ;
        RECT 1291.310 59.360 1291.590 59.640 ;
      LAYER met3 ;
        RECT 536.630 492.130 537.010 492.140 ;
        RECT 537.345 492.130 537.675 492.145 ;
        RECT 536.630 491.830 537.675 492.130 ;
        RECT 536.630 491.820 537.010 491.830 ;
        RECT 537.345 491.815 537.675 491.830 ;
        RECT 536.630 59.650 537.010 59.660 ;
        RECT 1291.285 59.650 1291.615 59.665 ;
        RECT 536.630 59.350 1291.615 59.650 ;
        RECT 536.630 59.340 537.010 59.350 ;
        RECT 1291.285 59.335 1291.615 59.350 ;
      LAYER via3 ;
        RECT 536.660 491.820 536.980 492.140 ;
        RECT 536.660 59.340 536.980 59.660 ;
      LAYER met4 ;
        RECT 536.655 491.815 536.985 492.145 ;
        RECT 536.670 59.665 536.970 491.815 ;
        RECT 536.655 59.335 536.985 59.665 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.040 499.500 538.360 499.760 ;
        RECT 538.130 498.400 538.270 499.500 ;
        RECT 538.130 498.200 538.590 498.400 ;
        RECT 538.270 498.140 538.590 498.200 ;
        RECT 538.270 51.920 538.590 51.980 ;
        RECT 1308.770 51.920 1309.090 51.980 ;
        RECT 538.270 51.780 1309.090 51.920 ;
        RECT 538.270 51.720 538.590 51.780 ;
        RECT 1308.770 51.720 1309.090 51.780 ;
      LAYER via ;
        RECT 538.070 499.500 538.330 499.760 ;
        RECT 538.300 498.140 538.560 498.400 ;
        RECT 538.300 51.720 538.560 51.980 ;
        RECT 1308.800 51.720 1309.060 51.980 ;
      LAYER met2 ;
        RECT 538.090 500.000 538.370 504.000 ;
        RECT 538.130 499.790 538.270 500.000 ;
        RECT 538.070 499.470 538.330 499.790 ;
        RECT 538.300 498.110 538.560 498.430 ;
        RECT 538.360 52.010 538.500 498.110 ;
        RECT 538.300 51.690 538.560 52.010 ;
        RECT 1308.800 51.690 1309.060 52.010 ;
        RECT 1308.860 2.400 1309.000 51.690 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 539.420 499.500 539.740 499.760 ;
        RECT 539.510 498.680 539.650 499.500 ;
        RECT 539.510 498.540 539.880 498.680 ;
        RECT 538.730 497.320 539.050 497.380 ;
        RECT 539.740 497.320 539.880 498.540 ;
        RECT 538.730 497.180 539.880 497.320 ;
        RECT 538.730 497.120 539.050 497.180 ;
        RECT 538.730 59.740 539.050 59.800 ;
        RECT 1324.870 59.740 1325.190 59.800 ;
        RECT 538.730 59.600 1325.190 59.740 ;
        RECT 538.730 59.540 539.050 59.600 ;
        RECT 1324.870 59.540 1325.190 59.600 ;
      LAYER via ;
        RECT 539.450 499.500 539.710 499.760 ;
        RECT 538.760 497.120 539.020 497.380 ;
        RECT 538.760 59.540 539.020 59.800 ;
        RECT 1324.900 59.540 1325.160 59.800 ;
      LAYER met2 ;
        RECT 539.470 500.000 539.750 504.000 ;
        RECT 539.510 499.790 539.650 500.000 ;
        RECT 539.450 499.470 539.710 499.790 ;
        RECT 538.760 497.090 539.020 497.410 ;
        RECT 538.820 59.830 538.960 497.090 ;
        RECT 538.760 59.510 539.020 59.830 ;
        RECT 1324.900 59.510 1325.160 59.830 ;
        RECT 1324.960 1.770 1325.100 59.510 ;
        RECT 1326.590 1.770 1327.150 2.400 ;
        RECT 1324.960 1.630 1327.150 1.770 ;
        RECT 1326.590 -4.800 1327.150 1.630 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 489.510 482.360 489.830 482.420 ;
        RECT 491.350 482.360 491.670 482.420 ;
        RECT 489.510 482.220 491.670 482.360 ;
        RECT 489.510 482.160 489.830 482.220 ;
        RECT 491.350 482.160 491.670 482.220 ;
        RECT 490.890 75.040 491.210 75.100 ;
        RECT 685.930 75.040 686.250 75.100 ;
        RECT 490.890 74.900 686.250 75.040 ;
        RECT 490.890 74.840 491.210 74.900 ;
        RECT 685.930 74.840 686.250 74.900 ;
      LAYER via ;
        RECT 489.540 482.160 489.800 482.420 ;
        RECT 491.380 482.160 491.640 482.420 ;
        RECT 490.920 74.840 491.180 75.100 ;
        RECT 685.960 74.840 686.220 75.100 ;
      LAYER met2 ;
        RECT 489.790 500.000 490.070 504.000 ;
        RECT 489.830 498.340 489.970 500.000 ;
        RECT 489.600 498.200 489.970 498.340 ;
        RECT 489.600 482.450 489.740 498.200 ;
        RECT 489.540 482.130 489.800 482.450 ;
        RECT 491.380 482.130 491.640 482.450 ;
        RECT 491.440 473.010 491.580 482.130 ;
        RECT 490.980 472.870 491.580 473.010 ;
        RECT 490.980 75.130 491.120 472.870 ;
        RECT 490.920 74.810 491.180 75.130 ;
        RECT 685.960 74.810 686.220 75.130 ;
        RECT 686.020 1.770 686.160 74.810 ;
        RECT 688.110 1.770 688.670 2.400 ;
        RECT 686.020 1.630 688.670 1.770 ;
        RECT 688.110 -4.800 688.670 1.630 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 539.190 59.400 539.510 59.460 ;
        RECT 1341.890 59.400 1342.210 59.460 ;
        RECT 539.190 59.260 1342.210 59.400 ;
        RECT 539.190 59.200 539.510 59.260 ;
        RECT 1341.890 59.200 1342.210 59.260 ;
      LAYER via ;
        RECT 539.220 59.200 539.480 59.460 ;
        RECT 1341.920 59.200 1342.180 59.460 ;
      LAYER met2 ;
        RECT 540.850 500.000 541.130 504.000 ;
        RECT 540.890 498.680 541.030 500.000 ;
        RECT 540.660 498.540 541.030 498.680 ;
        RECT 540.660 472.445 540.800 498.540 ;
        RECT 539.210 472.075 539.490 472.445 ;
        RECT 540.590 472.075 540.870 472.445 ;
        RECT 539.280 59.490 539.420 472.075 ;
        RECT 539.220 59.170 539.480 59.490 ;
        RECT 1341.920 59.170 1342.180 59.490 ;
        RECT 1341.980 1.770 1342.120 59.170 ;
        RECT 1344.070 1.770 1344.630 2.400 ;
        RECT 1341.980 1.630 1344.630 1.770 ;
        RECT 1344.070 -4.800 1344.630 1.630 ;
      LAYER via2 ;
        RECT 539.210 472.120 539.490 472.400 ;
        RECT 540.590 472.120 540.870 472.400 ;
      LAYER met3 ;
        RECT 539.185 472.410 539.515 472.425 ;
        RECT 540.565 472.410 540.895 472.425 ;
        RECT 539.185 472.110 540.895 472.410 ;
        RECT 539.185 472.095 539.515 472.110 ;
        RECT 540.565 472.095 540.895 472.110 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 542.180 499.700 542.500 499.760 ;
        RECT 541.350 499.560 542.500 499.700 ;
        RECT 541.350 497.320 541.490 499.560 ;
        RECT 542.180 499.500 542.500 499.560 ;
        RECT 542.410 497.320 542.730 497.380 ;
        RECT 541.350 497.180 542.730 497.320 ;
        RECT 542.410 497.120 542.730 497.180 ;
        RECT 541.490 481.000 541.810 481.060 ;
        RECT 542.410 481.000 542.730 481.060 ;
        RECT 541.490 480.860 542.730 481.000 ;
        RECT 541.490 480.800 541.810 480.860 ;
        RECT 542.410 480.800 542.730 480.860 ;
        RECT 539.650 471.480 539.970 471.540 ;
        RECT 541.490 471.480 541.810 471.540 ;
        RECT 539.650 471.340 541.810 471.480 ;
        RECT 539.650 471.280 539.970 471.340 ;
        RECT 541.490 471.280 541.810 471.340 ;
        RECT 539.650 59.060 539.970 59.120 ;
        RECT 1362.130 59.060 1362.450 59.120 ;
        RECT 539.650 58.920 1362.450 59.060 ;
        RECT 539.650 58.860 539.970 58.920 ;
        RECT 1362.130 58.860 1362.450 58.920 ;
      LAYER via ;
        RECT 542.210 499.500 542.470 499.760 ;
        RECT 542.440 497.120 542.700 497.380 ;
        RECT 541.520 480.800 541.780 481.060 ;
        RECT 542.440 480.800 542.700 481.060 ;
        RECT 539.680 471.280 539.940 471.540 ;
        RECT 541.520 471.280 541.780 471.540 ;
        RECT 539.680 58.860 539.940 59.120 ;
        RECT 1362.160 58.860 1362.420 59.120 ;
      LAYER met2 ;
        RECT 542.230 500.000 542.510 504.000 ;
        RECT 542.270 499.790 542.410 500.000 ;
        RECT 542.210 499.470 542.470 499.790 ;
        RECT 542.440 497.090 542.700 497.410 ;
        RECT 542.500 481.090 542.640 497.090 ;
        RECT 541.520 480.770 541.780 481.090 ;
        RECT 542.440 480.770 542.700 481.090 ;
        RECT 541.580 471.570 541.720 480.770 ;
        RECT 539.680 471.250 539.940 471.570 ;
        RECT 541.520 471.250 541.780 471.570 ;
        RECT 539.740 59.150 539.880 471.250 ;
        RECT 539.680 58.830 539.940 59.150 ;
        RECT 1362.160 58.830 1362.420 59.150 ;
        RECT 1362.220 2.400 1362.360 58.830 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.610 500.000 543.890 504.000 ;
        RECT 543.650 499.815 543.790 500.000 ;
        RECT 543.580 499.445 543.860 499.815 ;
        RECT 1380.550 58.635 1380.830 59.005 ;
        RECT 1380.620 17.410 1380.760 58.635 ;
        RECT 1380.160 17.270 1380.760 17.410 ;
        RECT 1380.160 2.400 1380.300 17.270 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
      LAYER via2 ;
        RECT 543.580 499.490 543.860 499.770 ;
        RECT 1380.550 58.680 1380.830 58.960 ;
      LAYER met3 ;
        RECT 542.150 499.610 542.530 499.620 ;
        RECT 543.555 499.610 543.885 499.795 ;
        RECT 542.150 499.465 543.885 499.610 ;
        RECT 542.150 499.310 543.870 499.465 ;
        RECT 542.150 499.300 542.530 499.310 ;
        RECT 543.070 58.970 543.450 58.980 ;
        RECT 1380.525 58.970 1380.855 58.985 ;
        RECT 543.070 58.670 1380.855 58.970 ;
        RECT 543.070 58.660 543.450 58.670 ;
        RECT 1380.525 58.655 1380.855 58.670 ;
      LAYER via3 ;
        RECT 542.180 499.300 542.500 499.620 ;
        RECT 543.100 58.660 543.420 58.980 ;
      LAYER met4 ;
        RECT 542.175 499.610 542.505 499.625 ;
        RECT 542.175 499.310 543.410 499.610 ;
        RECT 542.175 499.295 542.505 499.310 ;
        RECT 543.110 58.985 543.410 499.310 ;
        RECT 543.095 58.655 543.425 58.985 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.170 472.500 545.490 472.560 ;
        RECT 547.930 472.500 548.250 472.560 ;
        RECT 545.170 472.360 548.250 472.500 ;
        RECT 545.170 472.300 545.490 472.360 ;
        RECT 547.930 472.300 548.250 472.360 ;
        RECT 547.930 130.120 548.250 130.180 ;
        RECT 1393.870 130.120 1394.190 130.180 ;
        RECT 547.930 129.980 1394.190 130.120 ;
        RECT 547.930 129.920 548.250 129.980 ;
        RECT 1393.870 129.920 1394.190 129.980 ;
      LAYER via ;
        RECT 545.200 472.300 545.460 472.560 ;
        RECT 547.960 472.300 548.220 472.560 ;
        RECT 547.960 129.920 548.220 130.180 ;
        RECT 1393.900 129.920 1394.160 130.180 ;
      LAYER met2 ;
        RECT 544.990 500.000 545.270 504.000 ;
        RECT 545.030 498.680 545.170 500.000 ;
        RECT 544.800 498.540 545.170 498.680 ;
        RECT 544.800 483.070 544.940 498.540 ;
        RECT 544.800 482.930 545.400 483.070 ;
        RECT 545.260 472.590 545.400 482.930 ;
        RECT 545.200 472.270 545.460 472.590 ;
        RECT 547.960 472.270 548.220 472.590 ;
        RECT 548.020 130.210 548.160 472.270 ;
        RECT 547.960 129.890 548.220 130.210 ;
        RECT 1393.900 129.890 1394.160 130.210 ;
        RECT 1393.960 82.870 1394.100 129.890 ;
        RECT 1393.960 82.730 1395.480 82.870 ;
        RECT 1395.340 1.770 1395.480 82.730 ;
        RECT 1397.430 1.770 1397.990 2.400 ;
        RECT 1395.340 1.630 1397.990 1.770 ;
        RECT 1397.430 -4.800 1397.990 1.630 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 546.320 499.700 546.640 499.760 ;
        RECT 546.320 499.500 546.780 499.700 ;
        RECT 546.640 499.080 546.780 499.500 ;
        RECT 546.550 498.820 546.870 499.080 ;
        RECT 546.550 491.540 546.870 491.600 ;
        RECT 564.030 491.540 564.350 491.600 ;
        RECT 546.550 491.400 564.350 491.540 ;
        RECT 546.550 491.340 546.870 491.400 ;
        RECT 564.030 491.340 564.350 491.400 ;
        RECT 563.570 129.780 563.890 129.840 ;
        RECT 1414.570 129.780 1414.890 129.840 ;
        RECT 563.570 129.640 1414.890 129.780 ;
        RECT 563.570 129.580 563.890 129.640 ;
        RECT 1414.570 129.580 1414.890 129.640 ;
      LAYER via ;
        RECT 546.350 499.500 546.610 499.760 ;
        RECT 546.580 498.820 546.840 499.080 ;
        RECT 546.580 491.340 546.840 491.600 ;
        RECT 564.060 491.340 564.320 491.600 ;
        RECT 563.600 129.580 563.860 129.840 ;
        RECT 1414.600 129.580 1414.860 129.840 ;
      LAYER met2 ;
        RECT 546.370 500.000 546.650 504.000 ;
        RECT 546.410 499.790 546.550 500.000 ;
        RECT 546.350 499.470 546.610 499.790 ;
        RECT 546.580 498.790 546.840 499.110 ;
        RECT 546.640 491.630 546.780 498.790 ;
        RECT 546.580 491.310 546.840 491.630 ;
        RECT 564.060 491.310 564.320 491.630 ;
        RECT 564.120 476.170 564.260 491.310 ;
        RECT 563.660 476.030 564.260 476.170 ;
        RECT 563.660 129.870 563.800 476.030 ;
        RECT 563.600 129.550 563.860 129.870 ;
        RECT 1414.600 129.550 1414.860 129.870 ;
        RECT 1414.660 82.870 1414.800 129.550 ;
        RECT 1414.660 82.730 1415.720 82.870 ;
        RECT 1415.580 2.400 1415.720 82.730 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 548.850 129.440 549.170 129.500 ;
        RECT 1428.370 129.440 1428.690 129.500 ;
        RECT 548.850 129.300 1428.690 129.440 ;
        RECT 548.850 129.240 549.170 129.300 ;
        RECT 1428.370 129.240 1428.690 129.300 ;
      LAYER via ;
        RECT 548.880 129.240 549.140 129.500 ;
        RECT 1428.400 129.240 1428.660 129.500 ;
      LAYER met2 ;
        RECT 547.750 500.000 548.030 504.000 ;
        RECT 547.790 499.475 547.930 500.000 ;
        RECT 547.720 499.105 548.000 499.475 ;
        RECT 548.870 497.915 549.150 498.285 ;
        RECT 548.940 129.530 549.080 497.915 ;
        RECT 548.880 129.210 549.140 129.530 ;
        RECT 1428.400 129.210 1428.660 129.530 ;
        RECT 1428.460 82.870 1428.600 129.210 ;
        RECT 1428.460 82.730 1433.200 82.870 ;
        RECT 1433.060 2.400 1433.200 82.730 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
      LAYER via2 ;
        RECT 547.720 499.150 548.000 499.430 ;
        RECT 548.870 497.960 549.150 498.240 ;
      LAYER met3 ;
        RECT 547.695 499.125 548.025 499.455 ;
        RECT 547.710 498.250 548.010 499.125 ;
        RECT 548.845 498.250 549.175 498.265 ;
        RECT 547.710 497.950 549.175 498.250 ;
        RECT 548.845 497.935 549.175 497.950 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 549.080 499.500 549.400 499.760 ;
        RECT 548.390 497.660 548.710 497.720 ;
        RECT 549.170 497.660 549.310 499.500 ;
        RECT 548.390 497.520 549.310 497.660 ;
        RECT 548.390 497.460 548.710 497.520 ;
        RECT 548.390 129.100 548.710 129.160 ;
        RECT 1449.070 129.100 1449.390 129.160 ;
        RECT 548.390 128.960 1449.390 129.100 ;
        RECT 548.390 128.900 548.710 128.960 ;
        RECT 1449.070 128.900 1449.390 128.960 ;
      LAYER via ;
        RECT 549.110 499.500 549.370 499.760 ;
        RECT 548.420 497.460 548.680 497.720 ;
        RECT 548.420 128.900 548.680 129.160 ;
        RECT 1449.100 128.900 1449.360 129.160 ;
      LAYER met2 ;
        RECT 549.130 500.000 549.410 504.000 ;
        RECT 549.170 499.790 549.310 500.000 ;
        RECT 549.110 499.470 549.370 499.790 ;
        RECT 548.420 497.430 548.680 497.750 ;
        RECT 548.480 129.190 548.620 497.430 ;
        RECT 548.420 128.870 548.680 129.190 ;
        RECT 1449.100 128.870 1449.360 129.190 ;
        RECT 1449.160 1.770 1449.300 128.870 ;
        RECT 1450.790 1.770 1451.350 2.400 ;
        RECT 1449.160 1.630 1451.350 1.770 ;
        RECT 1450.790 -4.800 1451.350 1.630 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.170 471.820 545.490 471.880 ;
        RECT 549.310 471.820 549.630 471.880 ;
        RECT 545.170 471.680 549.630 471.820 ;
        RECT 545.170 471.620 545.490 471.680 ;
        RECT 549.310 471.620 549.630 471.680 ;
        RECT 545.170 67.900 545.490 67.960 ;
        RECT 1466.090 67.900 1466.410 67.960 ;
        RECT 545.170 67.760 1466.410 67.900 ;
        RECT 545.170 67.700 545.490 67.760 ;
        RECT 1466.090 67.700 1466.410 67.760 ;
      LAYER via ;
        RECT 545.200 471.620 545.460 471.880 ;
        RECT 549.340 471.620 549.600 471.880 ;
        RECT 545.200 67.700 545.460 67.960 ;
        RECT 1466.120 67.700 1466.380 67.960 ;
      LAYER met2 ;
        RECT 550.510 500.000 550.790 504.000 ;
        RECT 550.550 499.645 550.690 500.000 ;
        RECT 550.480 499.275 550.760 499.645 ;
        RECT 549.790 498.850 550.070 498.965 ;
        RECT 549.400 498.710 550.070 498.850 ;
        RECT 549.400 471.910 549.540 498.710 ;
        RECT 549.790 498.595 550.070 498.710 ;
        RECT 545.200 471.590 545.460 471.910 ;
        RECT 549.340 471.590 549.600 471.910 ;
        RECT 545.260 67.990 545.400 471.590 ;
        RECT 545.200 67.670 545.460 67.990 ;
        RECT 1466.120 67.670 1466.380 67.990 ;
        RECT 1466.180 1.770 1466.320 67.670 ;
        RECT 1468.270 1.770 1468.830 2.400 ;
        RECT 1466.180 1.630 1468.830 1.770 ;
        RECT 1468.270 -4.800 1468.830 1.630 ;
      LAYER via2 ;
        RECT 550.480 499.320 550.760 499.600 ;
        RECT 549.790 498.640 550.070 498.920 ;
      LAYER met3 ;
        RECT 550.455 499.295 550.785 499.625 ;
        RECT 549.765 498.930 550.095 498.945 ;
        RECT 550.470 498.930 550.770 499.295 ;
        RECT 549.765 498.630 550.770 498.930 ;
        RECT 549.765 498.615 550.095 498.630 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 551.840 499.360 552.160 499.420 ;
        RECT 551.700 499.160 552.160 499.360 ;
        RECT 551.700 498.340 551.840 499.160 ;
        RECT 552.530 498.340 552.850 498.400 ;
        RECT 551.700 498.200 552.850 498.340 ;
        RECT 552.530 498.140 552.850 498.200 ;
        RECT 552.530 67.560 552.850 67.620 ;
        RECT 1486.330 67.560 1486.650 67.620 ;
        RECT 552.530 67.420 1486.650 67.560 ;
        RECT 552.530 67.360 552.850 67.420 ;
        RECT 1486.330 67.360 1486.650 67.420 ;
      LAYER via ;
        RECT 551.870 499.160 552.130 499.420 ;
        RECT 552.560 498.140 552.820 498.400 ;
        RECT 552.560 67.360 552.820 67.620 ;
        RECT 1486.360 67.360 1486.620 67.620 ;
      LAYER met2 ;
        RECT 551.890 500.000 552.170 504.000 ;
        RECT 551.930 499.450 552.070 500.000 ;
        RECT 551.870 499.130 552.130 499.450 ;
        RECT 552.560 498.110 552.820 498.430 ;
        RECT 552.620 67.650 552.760 498.110 ;
        RECT 552.560 67.330 552.820 67.650 ;
        RECT 1486.360 67.330 1486.620 67.650 ;
        RECT 1486.420 2.400 1486.560 67.330 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 553.220 499.700 553.540 499.760 ;
        RECT 553.220 499.500 553.680 499.700 ;
        RECT 553.540 498.740 553.680 499.500 ;
        RECT 553.450 498.480 553.770 498.740 ;
        RECT 552.070 472.840 552.390 472.900 ;
        RECT 552.990 472.840 553.310 472.900 ;
        RECT 552.070 472.700 553.310 472.840 ;
        RECT 552.070 472.640 552.390 472.700 ;
        RECT 552.990 472.640 553.310 472.700 ;
        RECT 552.070 66.880 552.390 66.940 ;
        RECT 1497.830 66.880 1498.150 66.940 ;
        RECT 552.070 66.740 1498.150 66.880 ;
        RECT 552.070 66.680 552.390 66.740 ;
        RECT 1497.830 66.680 1498.150 66.740 ;
        RECT 1497.830 19.280 1498.150 19.340 ;
        RECT 1503.810 19.280 1504.130 19.340 ;
        RECT 1497.830 19.140 1504.130 19.280 ;
        RECT 1497.830 19.080 1498.150 19.140 ;
        RECT 1503.810 19.080 1504.130 19.140 ;
      LAYER via ;
        RECT 553.250 499.500 553.510 499.760 ;
        RECT 553.480 498.480 553.740 498.740 ;
        RECT 552.100 472.640 552.360 472.900 ;
        RECT 553.020 472.640 553.280 472.900 ;
        RECT 552.100 66.680 552.360 66.940 ;
        RECT 1497.860 66.680 1498.120 66.940 ;
        RECT 1497.860 19.080 1498.120 19.340 ;
        RECT 1503.840 19.080 1504.100 19.340 ;
      LAYER met2 ;
        RECT 553.270 500.000 553.550 504.000 ;
        RECT 553.310 499.790 553.450 500.000 ;
        RECT 553.250 499.470 553.510 499.790 ;
        RECT 553.480 498.450 553.740 498.770 ;
        RECT 553.540 491.540 553.680 498.450 ;
        RECT 553.080 491.400 553.680 491.540 ;
        RECT 553.080 472.930 553.220 491.400 ;
        RECT 552.100 472.610 552.360 472.930 ;
        RECT 553.020 472.610 553.280 472.930 ;
        RECT 552.160 66.970 552.300 472.610 ;
        RECT 552.100 66.650 552.360 66.970 ;
        RECT 1497.860 66.650 1498.120 66.970 ;
        RECT 1497.920 19.370 1498.060 66.650 ;
        RECT 1497.860 19.050 1498.120 19.370 ;
        RECT 1503.840 19.050 1504.100 19.370 ;
        RECT 1503.900 2.400 1504.040 19.050 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 492.270 147.800 492.590 147.860 ;
        RECT 703.870 147.800 704.190 147.860 ;
        RECT 492.270 147.660 704.190 147.800 ;
        RECT 492.270 147.600 492.590 147.660 ;
        RECT 703.870 147.600 704.190 147.660 ;
      LAYER via ;
        RECT 492.300 147.600 492.560 147.860 ;
        RECT 703.900 147.600 704.160 147.860 ;
      LAYER met2 ;
        RECT 491.170 500.000 491.450 504.000 ;
        RECT 491.210 499.700 491.350 500.000 ;
        RECT 491.210 499.645 491.580 499.700 ;
        RECT 491.210 499.560 491.650 499.645 ;
        RECT 491.370 499.275 491.650 499.560 ;
        RECT 492.290 497.915 492.570 498.285 ;
        RECT 492.360 147.890 492.500 497.915 ;
        RECT 492.300 147.570 492.560 147.890 ;
        RECT 703.900 147.570 704.160 147.890 ;
        RECT 703.960 82.870 704.100 147.570 ;
        RECT 703.960 82.730 706.400 82.870 ;
        RECT 706.260 2.400 706.400 82.730 ;
        RECT 706.050 -4.800 706.610 2.400 ;
      LAYER via2 ;
        RECT 491.370 499.320 491.650 499.600 ;
        RECT 492.290 497.960 492.570 498.240 ;
      LAYER met3 ;
        RECT 491.345 499.295 491.675 499.625 ;
        RECT 491.360 498.250 491.660 499.295 ;
        RECT 492.265 498.250 492.595 498.265 ;
        RECT 491.360 497.950 492.595 498.250 ;
        RECT 492.265 497.935 492.595 497.950 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 554.600 499.500 554.920 499.760 ;
        RECT 554.690 498.740 554.830 499.500 ;
        RECT 554.370 498.540 554.830 498.740 ;
        RECT 554.370 498.480 554.690 498.540 ;
        RECT 552.990 472.160 553.310 472.220 ;
        RECT 554.370 472.160 554.690 472.220 ;
        RECT 552.990 472.020 554.690 472.160 ;
        RECT 552.990 471.960 553.310 472.020 ;
        RECT 554.370 471.960 554.690 472.020 ;
        RECT 552.990 66.540 553.310 66.600 ;
        RECT 1519.450 66.540 1519.770 66.600 ;
        RECT 552.990 66.400 1519.770 66.540 ;
        RECT 552.990 66.340 553.310 66.400 ;
        RECT 1519.450 66.340 1519.770 66.400 ;
      LAYER via ;
        RECT 554.630 499.500 554.890 499.760 ;
        RECT 554.400 498.480 554.660 498.740 ;
        RECT 553.020 471.960 553.280 472.220 ;
        RECT 554.400 471.960 554.660 472.220 ;
        RECT 553.020 66.340 553.280 66.600 ;
        RECT 1519.480 66.340 1519.740 66.600 ;
      LAYER met2 ;
        RECT 554.650 500.000 554.930 504.000 ;
        RECT 554.690 499.790 554.830 500.000 ;
        RECT 554.630 499.470 554.890 499.790 ;
        RECT 554.400 498.450 554.660 498.770 ;
        RECT 554.460 472.250 554.600 498.450 ;
        RECT 553.020 471.930 553.280 472.250 ;
        RECT 554.400 471.930 554.660 472.250 ;
        RECT 553.080 66.630 553.220 471.930 ;
        RECT 553.020 66.310 553.280 66.630 ;
        RECT 1519.480 66.310 1519.740 66.630 ;
        RECT 1519.540 1.770 1519.680 66.310 ;
        RECT 1521.630 1.770 1522.190 2.400 ;
        RECT 1519.540 1.630 1522.190 1.770 ;
        RECT 1521.630 -4.800 1522.190 1.630 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 555.980 499.500 556.300 499.760 ;
        RECT 556.070 499.080 556.210 499.500 ;
        RECT 556.070 498.880 556.530 499.080 ;
        RECT 556.210 498.820 556.530 498.880 ;
        RECT 555.290 128.760 555.610 128.820 ;
        RECT 1538.770 128.760 1539.090 128.820 ;
        RECT 555.290 128.620 1539.090 128.760 ;
        RECT 555.290 128.560 555.610 128.620 ;
        RECT 1538.770 128.560 1539.090 128.620 ;
      LAYER via ;
        RECT 556.010 499.500 556.270 499.760 ;
        RECT 556.240 498.820 556.500 499.080 ;
        RECT 555.320 128.560 555.580 128.820 ;
        RECT 1538.800 128.560 1539.060 128.820 ;
      LAYER met2 ;
        RECT 556.030 500.000 556.310 504.000 ;
        RECT 556.070 499.790 556.210 500.000 ;
        RECT 556.010 499.470 556.270 499.790 ;
        RECT 556.240 498.790 556.500 499.110 ;
        RECT 556.300 483.070 556.440 498.790 ;
        RECT 555.840 482.930 556.440 483.070 ;
        RECT 555.840 476.170 555.980 482.930 ;
        RECT 555.380 476.030 555.980 476.170 ;
        RECT 555.380 128.850 555.520 476.030 ;
        RECT 555.320 128.530 555.580 128.850 ;
        RECT 1538.800 128.530 1539.060 128.850 ;
        RECT 1538.860 17.410 1539.000 128.530 ;
        RECT 1538.860 17.270 1539.920 17.410 ;
        RECT 1539.780 2.400 1539.920 17.270 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.410 500.000 557.690 504.000 ;
        RECT 557.450 499.815 557.590 500.000 ;
        RECT 557.380 499.445 557.660 499.815 ;
        RECT 1557.190 74.275 1557.470 74.645 ;
        RECT 1557.260 2.400 1557.400 74.275 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
      LAYER via2 ;
        RECT 557.380 499.490 557.660 499.770 ;
        RECT 1557.190 74.320 1557.470 74.600 ;
      LAYER met3 ;
        RECT 557.355 499.780 557.685 499.795 ;
        RECT 557.140 499.465 557.685 499.780 ;
        RECT 555.950 498.930 556.330 498.940 ;
        RECT 557.140 498.930 557.440 499.465 ;
        RECT 555.950 498.630 557.440 498.930 ;
        RECT 555.950 498.620 556.330 498.630 ;
        RECT 555.950 74.610 556.330 74.620 ;
        RECT 1557.165 74.610 1557.495 74.625 ;
        RECT 555.950 74.310 1557.495 74.610 ;
        RECT 555.950 74.300 556.330 74.310 ;
        RECT 1557.165 74.295 1557.495 74.310 ;
      LAYER via3 ;
        RECT 555.980 498.620 556.300 498.940 ;
        RECT 555.980 74.300 556.300 74.620 ;
      LAYER met4 ;
        RECT 555.975 498.615 556.305 498.945 ;
        RECT 555.990 74.625 556.290 498.615 ;
        RECT 555.975 74.295 556.305 74.625 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.740 499.500 559.060 499.760 ;
        RECT 558.830 498.740 558.970 499.500 ;
        RECT 558.830 498.540 559.290 498.740 ;
        RECT 558.970 498.480 559.290 498.540 ;
        RECT 558.970 472.160 559.290 472.220 ;
        RECT 560.810 472.160 561.130 472.220 ;
        RECT 558.970 472.020 561.130 472.160 ;
        RECT 558.970 471.960 559.290 472.020 ;
        RECT 560.810 471.960 561.130 472.020 ;
        RECT 560.810 150.520 561.130 150.580 ;
        RECT 1573.270 150.520 1573.590 150.580 ;
        RECT 560.810 150.380 1573.590 150.520 ;
        RECT 560.810 150.320 561.130 150.380 ;
        RECT 1573.270 150.320 1573.590 150.380 ;
      LAYER via ;
        RECT 558.770 499.500 559.030 499.760 ;
        RECT 559.000 498.480 559.260 498.740 ;
        RECT 559.000 471.960 559.260 472.220 ;
        RECT 560.840 471.960 561.100 472.220 ;
        RECT 560.840 150.320 561.100 150.580 ;
        RECT 1573.300 150.320 1573.560 150.580 ;
      LAYER met2 ;
        RECT 558.790 500.000 559.070 504.000 ;
        RECT 558.830 499.790 558.970 500.000 ;
        RECT 558.770 499.470 559.030 499.790 ;
        RECT 559.000 498.450 559.260 498.770 ;
        RECT 559.060 472.250 559.200 498.450 ;
        RECT 559.000 471.930 559.260 472.250 ;
        RECT 560.840 471.930 561.100 472.250 ;
        RECT 560.900 150.610 561.040 471.930 ;
        RECT 560.840 150.290 561.100 150.610 ;
        RECT 1573.300 150.290 1573.560 150.610 ;
        RECT 1573.360 1.770 1573.500 150.290 ;
        RECT 1574.990 1.770 1575.550 2.400 ;
        RECT 1573.360 1.630 1575.550 1.770 ;
        RECT 1574.990 -4.800 1575.550 1.630 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 560.120 499.700 560.440 499.760 ;
        RECT 560.120 499.560 560.810 499.700 ;
        RECT 560.120 499.500 560.440 499.560 ;
        RECT 560.670 498.740 560.810 499.560 ;
        RECT 560.350 498.540 560.810 498.740 ;
        RECT 560.350 498.480 560.670 498.540 ;
        RECT 561.270 150.180 561.590 150.240 ;
        RECT 1587.070 150.180 1587.390 150.240 ;
        RECT 561.270 150.040 1587.390 150.180 ;
        RECT 561.270 149.980 561.590 150.040 ;
        RECT 1587.070 149.980 1587.390 150.040 ;
      LAYER via ;
        RECT 560.150 499.500 560.410 499.760 ;
        RECT 560.380 498.480 560.640 498.740 ;
        RECT 561.300 149.980 561.560 150.240 ;
        RECT 1587.100 149.980 1587.360 150.240 ;
      LAYER met2 ;
        RECT 560.170 500.000 560.450 504.000 ;
        RECT 560.210 499.790 560.350 500.000 ;
        RECT 560.150 499.470 560.410 499.790 ;
        RECT 560.380 498.450 560.640 498.770 ;
        RECT 560.440 473.010 560.580 498.450 ;
        RECT 560.440 472.870 561.500 473.010 ;
        RECT 561.360 150.270 561.500 472.870 ;
        RECT 561.300 149.950 561.560 150.270 ;
        RECT 1587.100 149.950 1587.360 150.270 ;
        RECT 1587.160 82.870 1587.300 149.950 ;
        RECT 1587.160 82.730 1590.520 82.870 ;
        RECT 1590.380 1.770 1590.520 82.730 ;
        RECT 1592.470 1.770 1593.030 2.400 ;
        RECT 1590.380 1.630 1593.030 1.770 ;
        RECT 1592.470 -4.800 1593.030 1.630 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 561.500 499.360 561.820 499.420 ;
        RECT 561.500 499.160 561.960 499.360 ;
        RECT 561.820 498.400 561.960 499.160 ;
        RECT 561.730 498.140 562.050 498.400 ;
        RECT 561.730 474.000 562.050 474.260 ;
        RECT 559.430 471.820 559.750 471.880 ;
        RECT 561.820 471.820 561.960 474.000 ;
        RECT 559.430 471.680 561.960 471.820 ;
        RECT 559.430 471.620 559.750 471.680 ;
        RECT 559.430 66.200 559.750 66.260 ;
        RECT 1610.530 66.200 1610.850 66.260 ;
        RECT 559.430 66.060 1610.850 66.200 ;
        RECT 559.430 66.000 559.750 66.060 ;
        RECT 1610.530 66.000 1610.850 66.060 ;
      LAYER via ;
        RECT 561.530 499.160 561.790 499.420 ;
        RECT 561.760 498.140 562.020 498.400 ;
        RECT 561.760 474.000 562.020 474.260 ;
        RECT 559.460 471.620 559.720 471.880 ;
        RECT 559.460 66.000 559.720 66.260 ;
        RECT 1610.560 66.000 1610.820 66.260 ;
      LAYER met2 ;
        RECT 561.550 500.000 561.830 504.000 ;
        RECT 561.590 499.450 561.730 500.000 ;
        RECT 561.530 499.130 561.790 499.450 ;
        RECT 561.760 498.110 562.020 498.430 ;
        RECT 561.820 474.290 561.960 498.110 ;
        RECT 561.760 473.970 562.020 474.290 ;
        RECT 559.460 471.590 559.720 471.910 ;
        RECT 559.520 66.290 559.660 471.590 ;
        RECT 559.460 65.970 559.720 66.290 ;
        RECT 1610.560 65.970 1610.820 66.290 ;
        RECT 1610.620 2.400 1610.760 65.970 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 561.730 149.840 562.050 149.900 ;
        RECT 1621.570 149.840 1621.890 149.900 ;
        RECT 561.730 149.700 1621.890 149.840 ;
        RECT 561.730 149.640 562.050 149.700 ;
        RECT 1621.570 149.640 1621.890 149.700 ;
        RECT 1621.570 16.900 1621.890 16.960 ;
        RECT 1628.010 16.900 1628.330 16.960 ;
        RECT 1621.570 16.760 1628.330 16.900 ;
        RECT 1621.570 16.700 1621.890 16.760 ;
        RECT 1628.010 16.700 1628.330 16.760 ;
      LAYER via ;
        RECT 561.760 149.640 562.020 149.900 ;
        RECT 1621.600 149.640 1621.860 149.900 ;
        RECT 1621.600 16.700 1621.860 16.960 ;
        RECT 1628.040 16.700 1628.300 16.960 ;
      LAYER met2 ;
        RECT 562.930 500.000 563.210 504.000 ;
        RECT 562.970 498.170 563.110 500.000 ;
        RECT 562.970 498.030 563.340 498.170 ;
        RECT 563.200 476.170 563.340 498.030 ;
        RECT 562.740 476.030 563.340 476.170 ;
        RECT 562.740 470.970 562.880 476.030 ;
        RECT 561.820 470.830 562.880 470.970 ;
        RECT 561.820 149.930 561.960 470.830 ;
        RECT 561.760 149.610 562.020 149.930 ;
        RECT 1621.600 149.610 1621.860 149.930 ;
        RECT 1621.660 16.990 1621.800 149.610 ;
        RECT 1621.600 16.670 1621.860 16.990 ;
        RECT 1628.040 16.670 1628.300 16.990 ;
        RECT 1628.100 2.400 1628.240 16.670 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.310 500.000 564.590 504.000 ;
        RECT 564.350 499.815 564.490 500.000 ;
        RECT 564.280 499.445 564.560 499.815 ;
        RECT 1643.670 73.595 1643.950 73.965 ;
        RECT 1643.740 1.770 1643.880 73.595 ;
        RECT 1645.830 1.770 1646.390 2.400 ;
        RECT 1643.740 1.630 1646.390 1.770 ;
        RECT 1645.830 -4.800 1646.390 1.630 ;
      LAYER via2 ;
        RECT 564.280 499.490 564.560 499.770 ;
        RECT 1643.670 73.640 1643.950 73.920 ;
      LAYER met3 ;
        RECT 564.255 499.620 564.585 499.795 ;
        RECT 564.230 499.610 564.610 499.620 ;
        RECT 564.230 499.310 564.870 499.610 ;
        RECT 564.230 499.300 564.610 499.310 ;
        RECT 564.230 73.930 564.610 73.940 ;
        RECT 1643.645 73.930 1643.975 73.945 ;
        RECT 564.230 73.630 1643.975 73.930 ;
        RECT 564.230 73.620 564.610 73.630 ;
        RECT 1643.645 73.615 1643.975 73.630 ;
      LAYER via3 ;
        RECT 564.260 499.300 564.580 499.620 ;
        RECT 564.260 73.620 564.580 73.940 ;
      LAYER met4 ;
        RECT 564.255 499.295 564.585 499.625 ;
        RECT 564.270 73.945 564.570 499.295 ;
        RECT 564.255 73.615 564.585 73.945 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 565.870 497.660 566.190 497.720 ;
        RECT 568.170 497.660 568.490 497.720 ;
        RECT 565.870 497.520 568.490 497.660 ;
        RECT 565.870 497.460 566.190 497.520 ;
        RECT 568.170 497.460 568.490 497.520 ;
        RECT 566.790 472.840 567.110 472.900 ;
        RECT 568.170 472.840 568.490 472.900 ;
        RECT 566.790 472.700 568.490 472.840 ;
        RECT 566.790 472.640 567.110 472.700 ;
        RECT 568.170 472.640 568.490 472.700 ;
        RECT 566.790 73.680 567.110 73.740 ;
        RECT 1663.430 73.680 1663.750 73.740 ;
        RECT 566.790 73.540 1663.750 73.680 ;
        RECT 566.790 73.480 567.110 73.540 ;
        RECT 1663.430 73.480 1663.750 73.540 ;
      LAYER via ;
        RECT 565.900 497.460 566.160 497.720 ;
        RECT 568.200 497.460 568.460 497.720 ;
        RECT 566.820 472.640 567.080 472.900 ;
        RECT 568.200 472.640 568.460 472.900 ;
        RECT 566.820 73.480 567.080 73.740 ;
        RECT 1663.460 73.480 1663.720 73.740 ;
      LAYER met2 ;
        RECT 565.690 500.000 565.970 504.000 ;
        RECT 565.730 498.170 565.870 500.000 ;
        RECT 565.730 498.030 566.100 498.170 ;
        RECT 565.960 497.750 566.100 498.030 ;
        RECT 565.900 497.430 566.160 497.750 ;
        RECT 568.200 497.430 568.460 497.750 ;
        RECT 568.260 472.930 568.400 497.430 ;
        RECT 566.820 472.610 567.080 472.930 ;
        RECT 568.200 472.610 568.460 472.930 ;
        RECT 566.880 73.770 567.020 472.610 ;
        RECT 566.820 73.450 567.080 73.770 ;
        RECT 1663.460 73.450 1663.720 73.770 ;
        RECT 1663.520 2.400 1663.660 73.450 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 567.250 73.340 567.570 73.400 ;
        RECT 1681.370 73.340 1681.690 73.400 ;
        RECT 567.250 73.200 1681.690 73.340 ;
        RECT 567.250 73.140 567.570 73.200 ;
        RECT 1681.370 73.140 1681.690 73.200 ;
      LAYER via ;
        RECT 567.280 73.140 567.540 73.400 ;
        RECT 1681.400 73.140 1681.660 73.400 ;
      LAYER met2 ;
        RECT 567.070 500.000 567.350 504.000 ;
        RECT 567.110 499.645 567.250 500.000 ;
        RECT 567.040 499.275 567.320 499.645 ;
        RECT 566.810 497.915 567.090 498.285 ;
        RECT 566.880 492.050 567.020 497.915 ;
        RECT 566.880 491.910 567.480 492.050 ;
        RECT 567.340 73.430 567.480 491.910 ;
        RECT 567.280 73.110 567.540 73.430 ;
        RECT 1681.400 73.110 1681.660 73.430 ;
        RECT 1681.460 2.400 1681.600 73.110 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
      LAYER via2 ;
        RECT 567.040 499.320 567.320 499.600 ;
        RECT 566.810 497.960 567.090 498.240 ;
      LAYER met3 ;
        RECT 567.015 499.295 567.345 499.625 ;
        RECT 567.030 498.265 567.330 499.295 ;
        RECT 566.785 497.950 567.330 498.265 ;
        RECT 566.785 497.935 567.115 497.950 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 492.500 499.500 492.820 499.760 ;
        RECT 492.590 499.080 492.730 499.500 ;
        RECT 492.590 498.880 493.050 499.080 ;
        RECT 492.730 498.820 493.050 498.880 ;
        RECT 492.730 151.540 493.050 151.600 ;
        RECT 717.670 151.540 717.990 151.600 ;
        RECT 492.730 151.400 717.990 151.540 ;
        RECT 492.730 151.340 493.050 151.400 ;
        RECT 717.670 151.340 717.990 151.400 ;
        RECT 717.670 58.380 717.990 58.440 ;
        RECT 723.650 58.380 723.970 58.440 ;
        RECT 717.670 58.240 723.970 58.380 ;
        RECT 717.670 58.180 717.990 58.240 ;
        RECT 723.650 58.180 723.970 58.240 ;
      LAYER via ;
        RECT 492.530 499.500 492.790 499.760 ;
        RECT 492.760 498.820 493.020 499.080 ;
        RECT 492.760 151.340 493.020 151.600 ;
        RECT 717.700 151.340 717.960 151.600 ;
        RECT 717.700 58.180 717.960 58.440 ;
        RECT 723.680 58.180 723.940 58.440 ;
      LAYER met2 ;
        RECT 492.550 500.000 492.830 504.000 ;
        RECT 492.590 499.790 492.730 500.000 ;
        RECT 492.530 499.470 492.790 499.790 ;
        RECT 492.760 498.790 493.020 499.110 ;
        RECT 492.820 151.630 492.960 498.790 ;
        RECT 492.760 151.310 493.020 151.630 ;
        RECT 717.700 151.310 717.960 151.630 ;
        RECT 717.760 58.470 717.900 151.310 ;
        RECT 717.700 58.150 717.960 58.470 ;
        RECT 723.680 58.150 723.940 58.470 ;
        RECT 723.740 2.400 723.880 58.150 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.330 498.000 566.650 498.060 ;
        RECT 568.630 498.000 568.950 498.060 ;
        RECT 566.330 497.860 568.950 498.000 ;
        RECT 566.330 497.800 566.650 497.860 ;
        RECT 568.630 497.800 568.950 497.860 ;
        RECT 566.330 73.000 566.650 73.060 ;
        RECT 1697.470 73.000 1697.790 73.060 ;
        RECT 566.330 72.860 1697.790 73.000 ;
        RECT 566.330 72.800 566.650 72.860 ;
        RECT 1697.470 72.800 1697.790 72.860 ;
      LAYER via ;
        RECT 566.360 497.800 566.620 498.060 ;
        RECT 568.660 497.800 568.920 498.060 ;
        RECT 566.360 72.800 566.620 73.060 ;
        RECT 1697.500 72.800 1697.760 73.060 ;
      LAYER met2 ;
        RECT 568.450 500.000 568.730 504.000 ;
        RECT 568.490 498.680 568.630 500.000 ;
        RECT 568.490 498.540 568.860 498.680 ;
        RECT 568.720 498.090 568.860 498.540 ;
        RECT 566.360 497.770 566.620 498.090 ;
        RECT 568.660 497.770 568.920 498.090 ;
        RECT 566.420 73.090 566.560 497.770 ;
        RECT 566.360 72.770 566.620 73.090 ;
        RECT 1697.500 72.770 1697.760 73.090 ;
        RECT 1697.560 1.770 1697.700 72.770 ;
        RECT 1699.190 1.770 1699.750 2.400 ;
        RECT 1697.560 1.630 1699.750 1.770 ;
        RECT 1699.190 -4.800 1699.750 1.630 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 568.170 461.280 568.490 461.340 ;
        RECT 569.550 461.280 569.870 461.340 ;
        RECT 568.170 461.140 569.870 461.280 ;
        RECT 568.170 461.080 568.490 461.140 ;
        RECT 569.550 461.080 569.870 461.140 ;
        RECT 568.170 157.320 568.490 157.380 ;
        RECT 1711.270 157.320 1711.590 157.380 ;
        RECT 568.170 157.180 1711.590 157.320 ;
        RECT 568.170 157.120 568.490 157.180 ;
        RECT 1711.270 157.120 1711.590 157.180 ;
      LAYER via ;
        RECT 568.200 461.080 568.460 461.340 ;
        RECT 569.580 461.080 569.840 461.340 ;
        RECT 568.200 157.120 568.460 157.380 ;
        RECT 1711.300 157.120 1711.560 157.380 ;
      LAYER met2 ;
        RECT 569.830 500.000 570.110 504.000 ;
        RECT 569.870 499.815 570.010 500.000 ;
        RECT 569.800 499.445 570.080 499.815 ;
        RECT 569.570 497.915 569.850 498.285 ;
        RECT 569.640 461.370 569.780 497.915 ;
        RECT 568.200 461.050 568.460 461.370 ;
        RECT 569.580 461.050 569.840 461.370 ;
        RECT 568.260 157.410 568.400 461.050 ;
        RECT 568.200 157.090 568.460 157.410 ;
        RECT 1711.300 157.090 1711.560 157.410 ;
        RECT 1711.360 82.870 1711.500 157.090 ;
        RECT 1711.360 82.730 1714.720 82.870 ;
        RECT 1714.580 1.770 1714.720 82.730 ;
        RECT 1716.670 1.770 1717.230 2.400 ;
        RECT 1714.580 1.630 1717.230 1.770 ;
        RECT 1716.670 -4.800 1717.230 1.630 ;
      LAYER via2 ;
        RECT 569.800 499.490 570.080 499.770 ;
        RECT 569.570 497.960 569.850 498.240 ;
      LAYER met3 ;
        RECT 569.775 499.610 570.105 499.795 ;
        RECT 568.870 499.465 570.105 499.610 ;
        RECT 568.870 499.310 570.090 499.465 ;
        RECT 568.870 498.250 569.170 499.310 ;
        RECT 569.545 498.250 569.875 498.265 ;
        RECT 568.870 497.950 569.875 498.250 ;
        RECT 569.545 497.935 569.875 497.950 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 571.160 499.500 571.480 499.760 ;
        RECT 571.250 499.080 571.390 499.500 ;
        RECT 570.930 498.880 571.390 499.080 ;
        RECT 570.930 498.820 571.250 498.880 ;
      LAYER via ;
        RECT 571.190 499.500 571.450 499.760 ;
        RECT 570.960 498.820 571.220 499.080 ;
      LAYER met2 ;
        RECT 571.210 500.000 571.490 504.000 ;
        RECT 571.250 499.790 571.390 500.000 ;
        RECT 571.190 499.470 571.450 499.790 ;
        RECT 570.960 498.790 571.220 499.110 ;
        RECT 571.020 492.165 571.160 498.790 ;
        RECT 570.950 491.795 571.230 492.165 ;
        RECT 1734.750 81.755 1735.030 82.125 ;
        RECT 1734.820 2.400 1734.960 81.755 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
      LAYER via2 ;
        RECT 570.950 491.840 571.230 492.120 ;
        RECT 1734.750 81.800 1735.030 82.080 ;
      LAYER met3 ;
        RECT 568.830 492.130 569.210 492.140 ;
        RECT 570.925 492.130 571.255 492.145 ;
        RECT 568.830 491.830 571.255 492.130 ;
        RECT 568.830 491.820 569.210 491.830 ;
        RECT 570.925 491.815 571.255 491.830 ;
        RECT 568.830 82.090 569.210 82.100 ;
        RECT 1734.725 82.090 1735.055 82.105 ;
        RECT 568.830 81.790 1735.055 82.090 ;
        RECT 568.830 81.780 569.210 81.790 ;
        RECT 1734.725 81.775 1735.055 81.790 ;
      LAYER via3 ;
        RECT 568.860 491.820 569.180 492.140 ;
        RECT 568.860 81.780 569.180 82.100 ;
      LAYER met4 ;
        RECT 568.855 491.815 569.185 492.145 ;
        RECT 568.870 82.105 569.170 491.815 ;
        RECT 568.855 81.775 569.185 82.105 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 572.540 499.500 572.860 499.760 ;
        RECT 572.630 498.000 572.770 499.500 ;
        RECT 575.070 498.000 575.390 498.060 ;
        RECT 572.630 497.860 575.390 498.000 ;
        RECT 575.070 497.800 575.390 497.860 ;
        RECT 575.070 474.000 575.390 474.260 ;
        RECT 575.160 473.180 575.300 474.000 ;
        RECT 575.530 473.180 575.850 473.240 ;
        RECT 575.160 473.040 575.850 473.180 ;
        RECT 575.530 472.980 575.850 473.040 ;
        RECT 575.530 136.920 575.850 136.980 ;
        RECT 1745.770 136.920 1746.090 136.980 ;
        RECT 575.530 136.780 1746.090 136.920 ;
        RECT 575.530 136.720 575.850 136.780 ;
        RECT 1745.770 136.720 1746.090 136.780 ;
        RECT 1745.770 16.900 1746.090 16.960 ;
        RECT 1752.210 16.900 1752.530 16.960 ;
        RECT 1745.770 16.760 1752.530 16.900 ;
        RECT 1745.770 16.700 1746.090 16.760 ;
        RECT 1752.210 16.700 1752.530 16.760 ;
      LAYER via ;
        RECT 572.570 499.500 572.830 499.760 ;
        RECT 575.100 497.800 575.360 498.060 ;
        RECT 575.100 474.000 575.360 474.260 ;
        RECT 575.560 472.980 575.820 473.240 ;
        RECT 575.560 136.720 575.820 136.980 ;
        RECT 1745.800 136.720 1746.060 136.980 ;
        RECT 1745.800 16.700 1746.060 16.960 ;
        RECT 1752.240 16.700 1752.500 16.960 ;
      LAYER met2 ;
        RECT 572.590 500.000 572.870 504.000 ;
        RECT 572.630 499.790 572.770 500.000 ;
        RECT 572.570 499.470 572.830 499.790 ;
        RECT 575.100 497.770 575.360 498.090 ;
        RECT 575.160 474.290 575.300 497.770 ;
        RECT 575.100 473.970 575.360 474.290 ;
        RECT 575.560 472.950 575.820 473.270 ;
        RECT 575.620 137.010 575.760 472.950 ;
        RECT 575.560 136.690 575.820 137.010 ;
        RECT 1745.800 136.690 1746.060 137.010 ;
        RECT 1745.860 16.990 1746.000 136.690 ;
        RECT 1745.800 16.670 1746.060 16.990 ;
        RECT 1752.240 16.670 1752.500 16.990 ;
        RECT 1752.300 2.400 1752.440 16.670 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.150 472.840 574.470 472.900 ;
        RECT 576.450 472.840 576.770 472.900 ;
        RECT 574.150 472.700 576.770 472.840 ;
        RECT 574.150 472.640 574.470 472.700 ;
        RECT 576.450 472.640 576.770 472.700 ;
        RECT 576.450 156.980 576.770 157.040 ;
        RECT 1766.470 156.980 1766.790 157.040 ;
        RECT 576.450 156.840 1766.790 156.980 ;
        RECT 576.450 156.780 576.770 156.840 ;
        RECT 1766.470 156.780 1766.790 156.840 ;
      LAYER via ;
        RECT 574.180 472.640 574.440 472.900 ;
        RECT 576.480 472.640 576.740 472.900 ;
        RECT 576.480 156.780 576.740 157.040 ;
        RECT 1766.500 156.780 1766.760 157.040 ;
      LAYER met2 ;
        RECT 573.970 500.000 574.250 504.000 ;
        RECT 574.010 498.850 574.150 500.000 ;
        RECT 574.010 498.710 574.380 498.850 ;
        RECT 574.240 472.930 574.380 498.710 ;
        RECT 574.180 472.610 574.440 472.930 ;
        RECT 576.480 472.610 576.740 472.930 ;
        RECT 576.540 157.070 576.680 472.610 ;
        RECT 576.480 156.750 576.740 157.070 ;
        RECT 1766.500 156.750 1766.760 157.070 ;
        RECT 1766.560 82.870 1766.700 156.750 ;
        RECT 1766.560 82.730 1768.080 82.870 ;
        RECT 1767.940 1.770 1768.080 82.730 ;
        RECT 1770.030 1.770 1770.590 2.400 ;
        RECT 1767.940 1.630 1770.590 1.770 ;
        RECT 1770.030 -4.800 1770.590 1.630 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 573.230 80.480 573.550 80.540 ;
        RECT 1787.630 80.480 1787.950 80.540 ;
        RECT 573.230 80.340 1787.950 80.480 ;
        RECT 573.230 80.280 573.550 80.340 ;
        RECT 1787.630 80.280 1787.950 80.340 ;
      LAYER via ;
        RECT 573.260 80.280 573.520 80.540 ;
        RECT 1787.660 80.280 1787.920 80.540 ;
      LAYER met2 ;
        RECT 575.350 500.000 575.630 504.000 ;
        RECT 575.390 499.645 575.530 500.000 ;
        RECT 575.320 499.275 575.600 499.645 ;
        RECT 573.250 491.115 573.530 491.485 ;
        RECT 573.320 80.570 573.460 491.115 ;
        RECT 573.260 80.250 573.520 80.570 ;
        RECT 1787.660 80.250 1787.920 80.570 ;
        RECT 1787.720 2.400 1787.860 80.250 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
      LAYER via2 ;
        RECT 575.320 499.320 575.600 499.600 ;
        RECT 573.250 491.160 573.530 491.440 ;
      LAYER met3 ;
        RECT 575.295 499.620 575.625 499.625 ;
        RECT 575.270 499.610 575.650 499.620 ;
        RECT 575.270 499.310 576.080 499.610 ;
        RECT 575.270 499.300 575.650 499.310 ;
        RECT 575.295 499.295 575.625 499.300 ;
        RECT 573.225 491.450 573.555 491.465 ;
        RECT 575.270 491.450 575.650 491.460 ;
        RECT 573.225 491.150 575.650 491.450 ;
        RECT 573.225 491.135 573.555 491.150 ;
        RECT 575.270 491.140 575.650 491.150 ;
      LAYER via3 ;
        RECT 575.300 499.300 575.620 499.620 ;
        RECT 575.300 491.140 575.620 491.460 ;
      LAYER met4 ;
        RECT 575.295 499.295 575.625 499.625 ;
        RECT 575.310 491.465 575.610 499.295 ;
        RECT 575.295 491.135 575.625 491.465 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 576.680 499.360 577.000 499.420 ;
        RECT 576.080 499.220 577.000 499.360 ;
        RECT 576.080 498.400 576.220 499.220 ;
        RECT 576.680 499.160 577.000 499.220 ;
        RECT 575.990 498.140 576.310 498.400 ;
        RECT 575.990 156.640 576.310 156.700 ;
        RECT 1800.970 156.640 1801.290 156.700 ;
        RECT 575.990 156.500 1801.290 156.640 ;
        RECT 575.990 156.440 576.310 156.500 ;
        RECT 1800.970 156.440 1801.290 156.500 ;
      LAYER via ;
        RECT 576.710 499.160 576.970 499.420 ;
        RECT 576.020 498.140 576.280 498.400 ;
        RECT 576.020 156.440 576.280 156.700 ;
        RECT 1801.000 156.440 1801.260 156.700 ;
      LAYER met2 ;
        RECT 576.730 500.000 577.010 504.000 ;
        RECT 576.770 499.450 576.910 500.000 ;
        RECT 576.710 499.130 576.970 499.450 ;
        RECT 576.020 498.110 576.280 498.430 ;
        RECT 576.080 156.730 576.220 498.110 ;
        RECT 576.020 156.410 576.280 156.730 ;
        RECT 1801.000 156.410 1801.260 156.730 ;
        RECT 1801.060 82.870 1801.200 156.410 ;
        RECT 1801.060 82.730 1805.800 82.870 ;
        RECT 1805.660 2.400 1805.800 82.730 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.110 500.000 578.390 504.000 ;
        RECT 578.150 498.340 578.290 500.000 ;
        RECT 577.920 498.200 578.290 498.340 ;
        RECT 577.920 483.325 578.060 498.200 ;
        RECT 577.850 482.955 578.130 483.325 ;
        RECT 1823.070 81.075 1823.350 81.445 ;
        RECT 1823.140 2.400 1823.280 81.075 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
      LAYER via2 ;
        RECT 577.850 483.000 578.130 483.280 ;
        RECT 1823.070 81.120 1823.350 81.400 ;
      LAYER met3 ;
        RECT 577.825 483.300 578.155 483.305 ;
        RECT 577.825 483.290 578.410 483.300 ;
        RECT 577.600 482.990 578.410 483.290 ;
        RECT 577.825 482.980 578.410 482.990 ;
        RECT 577.825 482.975 578.155 482.980 ;
        RECT 578.030 81.410 578.410 81.420 ;
        RECT 1823.045 81.410 1823.375 81.425 ;
        RECT 578.030 81.110 1823.375 81.410 ;
        RECT 578.030 81.100 578.410 81.110 ;
        RECT 1823.045 81.095 1823.375 81.110 ;
      LAYER via3 ;
        RECT 578.060 482.980 578.380 483.300 ;
        RECT 578.060 81.100 578.380 81.420 ;
      LAYER met4 ;
        RECT 578.055 482.975 578.385 483.305 ;
        RECT 578.070 81.425 578.370 482.975 ;
        RECT 578.055 81.095 578.385 81.425 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 579.670 473.520 579.990 473.580 ;
        RECT 582.430 473.520 582.750 473.580 ;
        RECT 579.670 473.380 582.750 473.520 ;
        RECT 579.670 473.320 579.990 473.380 ;
        RECT 582.430 473.320 582.750 473.380 ;
        RECT 581.970 156.300 582.290 156.360 ;
        RECT 1835.470 156.300 1835.790 156.360 ;
        RECT 581.970 156.160 1835.790 156.300 ;
        RECT 581.970 156.100 582.290 156.160 ;
        RECT 1835.470 156.100 1835.790 156.160 ;
      LAYER via ;
        RECT 579.700 473.320 579.960 473.580 ;
        RECT 582.460 473.320 582.720 473.580 ;
        RECT 582.000 156.100 582.260 156.360 ;
        RECT 1835.500 156.100 1835.760 156.360 ;
      LAYER met2 ;
        RECT 579.490 500.000 579.770 504.000 ;
        RECT 579.530 498.680 579.670 500.000 ;
        RECT 579.530 498.540 579.900 498.680 ;
        RECT 579.760 473.610 579.900 498.540 ;
        RECT 579.700 473.290 579.960 473.610 ;
        RECT 582.460 473.290 582.720 473.610 ;
        RECT 582.520 472.330 582.660 473.290 ;
        RECT 582.060 472.190 582.660 472.330 ;
        RECT 582.060 156.390 582.200 472.190 ;
        RECT 582.000 156.070 582.260 156.390 ;
        RECT 1835.500 156.070 1835.760 156.390 ;
        RECT 1835.560 82.870 1835.700 156.070 ;
        RECT 1835.560 82.730 1838.920 82.870 ;
        RECT 1838.780 1.770 1838.920 82.730 ;
        RECT 1840.870 1.770 1841.430 2.400 ;
        RECT 1838.780 1.630 1841.430 1.770 ;
        RECT 1840.870 -4.800 1841.430 1.630 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 581.050 88.640 581.370 88.700 ;
        RECT 1856.170 88.640 1856.490 88.700 ;
        RECT 581.050 88.500 1856.490 88.640 ;
        RECT 581.050 88.440 581.370 88.500 ;
        RECT 1856.170 88.440 1856.490 88.500 ;
      LAYER via ;
        RECT 581.080 88.440 581.340 88.700 ;
        RECT 1856.200 88.440 1856.460 88.700 ;
      LAYER met2 ;
        RECT 580.870 500.000 581.150 504.000 ;
        RECT 580.910 499.700 581.050 500.000 ;
        RECT 580.910 499.560 581.280 499.700 ;
        RECT 581.140 88.730 581.280 499.560 ;
        RECT 581.080 88.410 581.340 88.730 ;
        RECT 1856.200 88.410 1856.460 88.730 ;
        RECT 1856.260 1.770 1856.400 88.410 ;
        RECT 1858.350 1.770 1858.910 2.400 ;
        RECT 1856.260 1.630 1858.910 1.770 ;
        RECT 1858.350 -4.800 1858.910 1.630 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 493.880 499.500 494.200 499.760 ;
        RECT 493.970 498.400 494.110 499.500 ;
        RECT 493.970 498.200 494.430 498.400 ;
        RECT 494.110 498.140 494.430 498.200 ;
        RECT 494.110 488.960 494.430 489.220 ;
        RECT 493.650 488.140 493.970 488.200 ;
        RECT 494.200 488.140 494.340 488.960 ;
        RECT 493.650 488.000 494.340 488.140 ;
        RECT 493.650 487.940 493.970 488.000 ;
        RECT 491.350 472.500 491.670 472.560 ;
        RECT 493.650 472.500 493.970 472.560 ;
        RECT 491.350 472.360 493.970 472.500 ;
        RECT 491.350 472.300 491.670 472.360 ;
        RECT 493.650 472.300 493.970 472.360 ;
        RECT 491.350 81.500 491.670 81.560 ;
        RECT 739.290 81.500 739.610 81.560 ;
        RECT 491.350 81.360 739.610 81.500 ;
        RECT 491.350 81.300 491.670 81.360 ;
        RECT 739.290 81.300 739.610 81.360 ;
      LAYER via ;
        RECT 493.910 499.500 494.170 499.760 ;
        RECT 494.140 498.140 494.400 498.400 ;
        RECT 494.140 488.960 494.400 489.220 ;
        RECT 493.680 487.940 493.940 488.200 ;
        RECT 491.380 472.300 491.640 472.560 ;
        RECT 493.680 472.300 493.940 472.560 ;
        RECT 491.380 81.300 491.640 81.560 ;
        RECT 739.320 81.300 739.580 81.560 ;
      LAYER met2 ;
        RECT 493.930 500.000 494.210 504.000 ;
        RECT 493.970 499.790 494.110 500.000 ;
        RECT 493.910 499.470 494.170 499.790 ;
        RECT 494.140 498.110 494.400 498.430 ;
        RECT 494.200 489.250 494.340 498.110 ;
        RECT 494.140 488.930 494.400 489.250 ;
        RECT 493.680 487.910 493.940 488.230 ;
        RECT 493.740 472.590 493.880 487.910 ;
        RECT 491.380 472.270 491.640 472.590 ;
        RECT 493.680 472.270 493.940 472.590 ;
        RECT 491.440 81.590 491.580 472.270 ;
        RECT 491.380 81.270 491.640 81.590 ;
        RECT 739.320 81.270 739.580 81.590 ;
        RECT 739.380 1.770 739.520 81.270 ;
        RECT 741.470 1.770 742.030 2.400 ;
        RECT 739.380 1.630 742.030 1.770 ;
        RECT 741.470 -4.800 742.030 1.630 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.590 472.840 580.910 472.900 ;
        RECT 581.970 472.840 582.290 472.900 ;
        RECT 580.590 472.700 582.290 472.840 ;
        RECT 580.590 472.640 580.910 472.700 ;
        RECT 581.970 472.640 582.290 472.700 ;
        RECT 580.590 88.300 580.910 88.360 ;
        RECT 1870.430 88.300 1870.750 88.360 ;
        RECT 580.590 88.160 1870.750 88.300 ;
        RECT 580.590 88.100 580.910 88.160 ;
        RECT 1870.430 88.100 1870.750 88.160 ;
        RECT 1870.430 16.900 1870.750 16.960 ;
        RECT 1876.410 16.900 1876.730 16.960 ;
        RECT 1870.430 16.760 1876.730 16.900 ;
        RECT 1870.430 16.700 1870.750 16.760 ;
        RECT 1876.410 16.700 1876.730 16.760 ;
      LAYER via ;
        RECT 580.620 472.640 580.880 472.900 ;
        RECT 582.000 472.640 582.260 472.900 ;
        RECT 580.620 88.100 580.880 88.360 ;
        RECT 1870.460 88.100 1870.720 88.360 ;
        RECT 1870.460 16.700 1870.720 16.960 ;
        RECT 1876.440 16.700 1876.700 16.960 ;
      LAYER met2 ;
        RECT 582.250 500.000 582.530 504.000 ;
        RECT 582.290 499.360 582.430 500.000 ;
        RECT 582.060 499.220 582.430 499.360 ;
        RECT 582.060 498.680 582.200 499.220 ;
        RECT 581.830 498.540 582.200 498.680 ;
        RECT 581.830 498.170 581.970 498.540 ;
        RECT 581.830 498.030 582.200 498.170 ;
        RECT 582.060 472.930 582.200 498.030 ;
        RECT 580.620 472.610 580.880 472.930 ;
        RECT 582.000 472.610 582.260 472.930 ;
        RECT 580.680 88.390 580.820 472.610 ;
        RECT 580.620 88.070 580.880 88.390 ;
        RECT 1870.460 88.070 1870.720 88.390 ;
        RECT 1870.520 16.990 1870.660 88.070 ;
        RECT 1870.460 16.670 1870.720 16.990 ;
        RECT 1876.440 16.670 1876.700 16.990 ;
        RECT 1876.500 2.400 1876.640 16.670 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 583.580 499.500 583.900 499.760 ;
        RECT 583.670 499.360 583.810 499.500 ;
        RECT 583.440 499.220 583.810 499.360 ;
        RECT 583.440 498.680 583.580 499.220 ;
        RECT 584.270 498.680 584.590 498.740 ;
        RECT 583.440 498.540 584.590 498.680 ;
        RECT 584.270 498.480 584.590 498.540 ;
        RECT 580.130 472.500 580.450 472.560 ;
        RECT 583.810 472.500 584.130 472.560 ;
        RECT 580.130 472.360 584.130 472.500 ;
        RECT 580.130 472.300 580.450 472.360 ;
        RECT 583.810 472.300 584.130 472.360 ;
        RECT 580.130 45.120 580.450 45.180 ;
        RECT 1894.350 45.120 1894.670 45.180 ;
        RECT 580.130 44.980 1894.670 45.120 ;
        RECT 580.130 44.920 580.450 44.980 ;
        RECT 1894.350 44.920 1894.670 44.980 ;
      LAYER via ;
        RECT 583.610 499.500 583.870 499.760 ;
        RECT 584.300 498.480 584.560 498.740 ;
        RECT 580.160 472.300 580.420 472.560 ;
        RECT 583.840 472.300 584.100 472.560 ;
        RECT 580.160 44.920 580.420 45.180 ;
        RECT 1894.380 44.920 1894.640 45.180 ;
      LAYER met2 ;
        RECT 583.630 500.000 583.910 504.000 ;
        RECT 583.670 499.790 583.810 500.000 ;
        RECT 583.610 499.470 583.870 499.790 ;
        RECT 584.300 498.450 584.560 498.770 ;
        RECT 584.360 490.010 584.500 498.450 ;
        RECT 583.900 489.870 584.500 490.010 ;
        RECT 583.900 472.590 584.040 489.870 ;
        RECT 580.160 472.270 580.420 472.590 ;
        RECT 583.840 472.270 584.100 472.590 ;
        RECT 580.220 45.210 580.360 472.270 ;
        RECT 580.160 44.890 580.420 45.210 ;
        RECT 1894.380 44.890 1894.640 45.210 ;
        RECT 1894.440 2.400 1894.580 44.890 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.010 500.000 585.290 504.000 ;
        RECT 585.050 499.645 585.190 500.000 ;
        RECT 584.980 499.275 585.260 499.645 ;
        RECT 1911.850 80.395 1912.130 80.765 ;
        RECT 1911.920 2.400 1912.060 80.395 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
      LAYER via2 ;
        RECT 584.980 499.320 585.260 499.600 ;
        RECT 1911.850 80.440 1912.130 80.720 ;
      LAYER met3 ;
        RECT 583.550 499.610 583.930 499.620 ;
        RECT 584.955 499.610 585.285 499.625 ;
        RECT 583.550 499.310 585.285 499.610 ;
        RECT 583.550 499.300 583.930 499.310 ;
        RECT 584.955 499.295 585.285 499.310 ;
        RECT 583.550 80.730 583.930 80.740 ;
        RECT 1911.825 80.730 1912.155 80.745 ;
        RECT 583.550 80.430 1912.155 80.730 ;
        RECT 583.550 80.420 583.930 80.430 ;
        RECT 1911.825 80.415 1912.155 80.430 ;
      LAYER via3 ;
        RECT 583.580 499.300 583.900 499.620 ;
        RECT 583.580 80.420 583.900 80.740 ;
      LAYER met4 ;
        RECT 583.575 499.295 583.905 499.625 ;
        RECT 583.590 80.745 583.890 499.295 ;
        RECT 583.575 80.415 583.905 80.745 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.340 499.500 586.660 499.760 ;
        RECT 586.430 499.080 586.570 499.500 ;
        RECT 586.430 498.880 586.890 499.080 ;
        RECT 586.570 498.820 586.890 498.880 ;
        RECT 586.570 87.960 586.890 88.020 ;
        RECT 1925.170 87.960 1925.490 88.020 ;
        RECT 586.570 87.820 1925.490 87.960 ;
        RECT 586.570 87.760 586.890 87.820 ;
        RECT 1925.170 87.760 1925.490 87.820 ;
      LAYER via ;
        RECT 586.370 499.500 586.630 499.760 ;
        RECT 586.600 498.820 586.860 499.080 ;
        RECT 586.600 87.760 586.860 88.020 ;
        RECT 1925.200 87.760 1925.460 88.020 ;
      LAYER met2 ;
        RECT 586.390 500.000 586.670 504.000 ;
        RECT 586.430 499.790 586.570 500.000 ;
        RECT 586.370 499.470 586.630 499.790 ;
        RECT 586.600 498.790 586.860 499.110 ;
        RECT 586.660 88.050 586.800 498.790 ;
        RECT 586.600 87.730 586.860 88.050 ;
        RECT 1925.200 87.730 1925.460 88.050 ;
        RECT 1925.260 82.870 1925.400 87.730 ;
        RECT 1925.260 82.730 1928.160 82.870 ;
        RECT 1928.020 17.410 1928.160 82.730 ;
        RECT 1928.020 17.270 1930.000 17.410 ;
        RECT 1929.860 2.400 1930.000 17.270 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 587.490 87.620 587.810 87.680 ;
        RECT 1945.870 87.620 1946.190 87.680 ;
        RECT 587.490 87.480 1946.190 87.620 ;
        RECT 587.490 87.420 587.810 87.480 ;
        RECT 1945.870 87.420 1946.190 87.480 ;
      LAYER via ;
        RECT 587.520 87.420 587.780 87.680 ;
        RECT 1945.900 87.420 1946.160 87.680 ;
      LAYER met2 ;
        RECT 587.770 500.000 588.050 504.000 ;
        RECT 587.810 499.815 587.950 500.000 ;
        RECT 587.740 499.445 588.020 499.815 ;
        RECT 587.510 497.915 587.790 498.285 ;
        RECT 587.580 87.710 587.720 497.915 ;
        RECT 587.520 87.390 587.780 87.710 ;
        RECT 1945.900 87.390 1946.160 87.710 ;
        RECT 1945.960 82.870 1946.100 87.390 ;
        RECT 1945.960 82.730 1947.480 82.870 ;
        RECT 1947.340 2.400 1947.480 82.730 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
      LAYER via2 ;
        RECT 587.740 499.490 588.020 499.770 ;
        RECT 587.510 497.960 587.790 498.240 ;
      LAYER met3 ;
        RECT 587.715 499.780 588.045 499.795 ;
        RECT 587.500 499.465 588.045 499.780 ;
        RECT 587.500 498.265 587.800 499.465 ;
        RECT 587.485 497.935 587.815 498.265 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 589.100 499.160 589.420 499.420 ;
        RECT 589.190 499.020 589.330 499.160 ;
        RECT 588.960 498.880 589.330 499.020 ;
        RECT 588.960 498.400 589.100 498.880 ;
        RECT 588.870 498.140 589.190 498.400 ;
        RECT 587.030 491.880 587.350 491.940 ;
        RECT 588.870 491.880 589.190 491.940 ;
        RECT 587.030 491.740 589.190 491.880 ;
        RECT 587.030 491.680 587.350 491.740 ;
        RECT 588.870 491.680 589.190 491.740 ;
        RECT 587.030 87.280 587.350 87.340 ;
        RECT 1959.670 87.280 1959.990 87.340 ;
        RECT 587.030 87.140 1959.990 87.280 ;
        RECT 587.030 87.080 587.350 87.140 ;
        RECT 1959.670 87.080 1959.990 87.140 ;
      LAYER via ;
        RECT 589.130 499.160 589.390 499.420 ;
        RECT 588.900 498.140 589.160 498.400 ;
        RECT 587.060 491.680 587.320 491.940 ;
        RECT 588.900 491.680 589.160 491.940 ;
        RECT 587.060 87.080 587.320 87.340 ;
        RECT 1959.700 87.080 1959.960 87.340 ;
      LAYER met2 ;
        RECT 589.150 500.000 589.430 504.000 ;
        RECT 589.190 499.450 589.330 500.000 ;
        RECT 589.130 499.130 589.390 499.450 ;
        RECT 588.900 498.110 589.160 498.430 ;
        RECT 588.960 491.970 589.100 498.110 ;
        RECT 587.060 491.650 587.320 491.970 ;
        RECT 588.900 491.650 589.160 491.970 ;
        RECT 587.120 87.370 587.260 491.650 ;
        RECT 587.060 87.050 587.320 87.370 ;
        RECT 1959.700 87.050 1959.960 87.370 ;
        RECT 1959.760 82.870 1959.900 87.050 ;
        RECT 1959.760 82.730 1963.120 82.870 ;
        RECT 1962.980 1.770 1963.120 82.730 ;
        RECT 1965.070 1.770 1965.630 2.400 ;
        RECT 1962.980 1.630 1965.630 1.770 ;
        RECT 1965.070 -4.800 1965.630 1.630 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 590.250 491.880 590.570 491.940 ;
        RECT 591.170 491.880 591.490 491.940 ;
        RECT 590.250 491.740 591.490 491.880 ;
        RECT 590.250 491.680 590.570 491.740 ;
        RECT 591.170 491.680 591.490 491.740 ;
        RECT 588.870 473.520 589.190 473.580 ;
        RECT 590.250 473.520 590.570 473.580 ;
        RECT 588.870 473.380 590.570 473.520 ;
        RECT 588.870 473.320 589.190 473.380 ;
        RECT 590.250 473.320 590.570 473.380 ;
        RECT 588.870 155.960 589.190 156.020 ;
        RECT 1980.370 155.960 1980.690 156.020 ;
        RECT 588.870 155.820 1980.690 155.960 ;
        RECT 588.870 155.760 589.190 155.820 ;
        RECT 1980.370 155.760 1980.690 155.820 ;
      LAYER via ;
        RECT 590.280 491.680 590.540 491.940 ;
        RECT 591.200 491.680 591.460 491.940 ;
        RECT 588.900 473.320 589.160 473.580 ;
        RECT 590.280 473.320 590.540 473.580 ;
        RECT 588.900 155.760 589.160 156.020 ;
        RECT 1980.400 155.760 1980.660 156.020 ;
      LAYER met2 ;
        RECT 590.530 500.000 590.810 504.000 ;
        RECT 590.570 499.020 590.710 500.000 ;
        RECT 590.340 498.880 590.710 499.020 ;
        RECT 590.340 498.285 590.480 498.880 ;
        RECT 590.270 497.915 590.550 498.285 ;
        RECT 591.190 497.915 591.470 498.285 ;
        RECT 591.260 491.970 591.400 497.915 ;
        RECT 590.280 491.650 590.540 491.970 ;
        RECT 591.200 491.650 591.460 491.970 ;
        RECT 590.340 473.610 590.480 491.650 ;
        RECT 588.900 473.290 589.160 473.610 ;
        RECT 590.280 473.290 590.540 473.610 ;
        RECT 588.960 156.050 589.100 473.290 ;
        RECT 588.900 155.730 589.160 156.050 ;
        RECT 1980.400 155.730 1980.660 156.050 ;
        RECT 1980.460 1.770 1980.600 155.730 ;
        RECT 1982.550 1.770 1983.110 2.400 ;
        RECT 1980.460 1.630 1983.110 1.770 ;
        RECT 1982.550 -4.800 1983.110 1.630 ;
      LAYER via2 ;
        RECT 590.270 497.960 590.550 498.240 ;
        RECT 591.190 497.960 591.470 498.240 ;
      LAYER met3 ;
        RECT 590.245 498.250 590.575 498.265 ;
        RECT 591.165 498.250 591.495 498.265 ;
        RECT 590.245 497.950 591.495 498.250 ;
        RECT 590.245 497.935 590.575 497.950 ;
        RECT 591.165 497.935 591.495 497.950 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1994.170 16.900 1994.490 16.960 ;
        RECT 2000.610 16.900 2000.930 16.960 ;
        RECT 1994.170 16.760 2000.930 16.900 ;
        RECT 1994.170 16.700 1994.490 16.760 ;
        RECT 2000.610 16.700 2000.930 16.760 ;
      LAYER via ;
        RECT 1994.200 16.700 1994.460 16.960 ;
        RECT 2000.640 16.700 2000.900 16.960 ;
      LAYER met2 ;
        RECT 591.910 500.000 592.190 504.000 ;
        RECT 591.950 498.850 592.090 500.000 ;
        RECT 591.030 498.710 592.090 498.850 ;
        RECT 591.030 498.680 591.170 498.710 ;
        RECT 590.800 498.540 591.170 498.680 ;
        RECT 590.800 493.525 590.940 498.540 ;
        RECT 590.730 493.155 591.010 493.525 ;
        RECT 1994.190 130.035 1994.470 130.405 ;
        RECT 1994.260 16.990 1994.400 130.035 ;
        RECT 1994.200 16.670 1994.460 16.990 ;
        RECT 2000.640 16.670 2000.900 16.990 ;
        RECT 2000.700 2.400 2000.840 16.670 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
      LAYER via2 ;
        RECT 590.730 493.200 591.010 493.480 ;
        RECT 1994.190 130.080 1994.470 130.360 ;
      LAYER met3 ;
        RECT 590.705 493.500 591.035 493.505 ;
        RECT 590.705 493.490 591.290 493.500 ;
        RECT 590.705 493.190 591.490 493.490 ;
        RECT 590.705 493.180 591.290 493.190 ;
        RECT 590.705 493.175 591.035 493.180 ;
        RECT 590.910 130.370 591.290 130.380 ;
        RECT 1994.165 130.370 1994.495 130.385 ;
        RECT 590.910 130.070 1994.495 130.370 ;
        RECT 590.910 130.060 591.290 130.070 ;
        RECT 1994.165 130.055 1994.495 130.070 ;
      LAYER via3 ;
        RECT 590.940 493.180 591.260 493.500 ;
        RECT 590.940 130.060 591.260 130.380 ;
      LAYER met4 ;
        RECT 590.935 493.175 591.265 493.505 ;
        RECT 590.950 130.385 591.250 493.175 ;
        RECT 590.935 130.055 591.265 130.385 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.240 499.500 593.560 499.760 ;
        RECT 593.330 498.680 593.470 499.500 ;
        RECT 593.330 498.540 593.930 498.680 ;
        RECT 593.790 497.040 593.930 498.540 ;
        RECT 593.790 496.840 594.250 497.040 ;
        RECT 593.930 496.780 594.250 496.840 ;
        RECT 593.930 472.160 594.250 472.220 ;
        RECT 596.690 472.160 597.010 472.220 ;
        RECT 593.930 472.020 597.010 472.160 ;
        RECT 593.930 471.960 594.250 472.020 ;
        RECT 596.690 471.960 597.010 472.020 ;
        RECT 596.690 163.100 597.010 163.160 ;
        RECT 2014.870 163.100 2015.190 163.160 ;
        RECT 596.690 162.960 2015.190 163.100 ;
        RECT 596.690 162.900 597.010 162.960 ;
        RECT 2014.870 162.900 2015.190 162.960 ;
      LAYER via ;
        RECT 593.270 499.500 593.530 499.760 ;
        RECT 593.960 496.780 594.220 497.040 ;
        RECT 593.960 471.960 594.220 472.220 ;
        RECT 596.720 471.960 596.980 472.220 ;
        RECT 596.720 162.900 596.980 163.160 ;
        RECT 2014.900 162.900 2015.160 163.160 ;
      LAYER met2 ;
        RECT 593.290 500.000 593.570 504.000 ;
        RECT 593.330 499.790 593.470 500.000 ;
        RECT 593.270 499.470 593.530 499.790 ;
        RECT 593.960 496.750 594.220 497.070 ;
        RECT 594.020 472.250 594.160 496.750 ;
        RECT 593.960 471.930 594.220 472.250 ;
        RECT 596.720 471.930 596.980 472.250 ;
        RECT 596.780 163.190 596.920 471.930 ;
        RECT 596.720 162.870 596.980 163.190 ;
        RECT 2014.900 162.870 2015.160 163.190 ;
        RECT 2014.960 82.870 2015.100 162.870 ;
        RECT 2014.960 82.730 2018.320 82.870 ;
        RECT 2018.180 2.400 2018.320 82.730 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.470 86.940 593.790 87.000 ;
        RECT 2036.030 86.940 2036.350 87.000 ;
        RECT 593.470 86.800 2036.350 86.940 ;
        RECT 593.470 86.740 593.790 86.800 ;
        RECT 2036.030 86.740 2036.350 86.800 ;
      LAYER via ;
        RECT 593.500 86.740 593.760 87.000 ;
        RECT 2036.060 86.740 2036.320 87.000 ;
      LAYER met2 ;
        RECT 594.670 500.000 594.950 504.000 ;
        RECT 594.710 499.815 594.850 500.000 ;
        RECT 594.640 499.445 594.920 499.815 ;
        RECT 593.490 498.595 593.770 498.965 ;
        RECT 593.560 87.030 593.700 498.595 ;
        RECT 593.500 86.710 593.760 87.030 ;
        RECT 2036.060 86.710 2036.320 87.030 ;
        RECT 2036.120 2.400 2036.260 86.710 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
      LAYER via2 ;
        RECT 594.640 499.490 594.920 499.770 ;
        RECT 593.490 498.640 593.770 498.920 ;
      LAYER met3 ;
        RECT 594.615 499.465 594.945 499.795 ;
        RECT 593.465 498.930 593.795 498.945 ;
        RECT 594.630 498.930 594.930 499.465 ;
        RECT 593.465 498.630 594.930 498.930 ;
        RECT 593.465 498.615 593.795 498.630 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 501.010 164.800 501.330 164.860 ;
        RECT 759.070 164.800 759.390 164.860 ;
        RECT 501.010 164.660 759.390 164.800 ;
        RECT 501.010 164.600 501.330 164.660 ;
        RECT 759.070 164.600 759.390 164.660 ;
      LAYER via ;
        RECT 501.040 164.600 501.300 164.860 ;
        RECT 759.100 164.600 759.360 164.860 ;
      LAYER met2 ;
        RECT 495.310 500.000 495.590 504.000 ;
        RECT 495.350 499.645 495.490 500.000 ;
        RECT 495.280 499.275 495.560 499.645 ;
        RECT 501.030 489.755 501.310 490.125 ;
        RECT 501.100 164.890 501.240 489.755 ;
        RECT 501.040 164.570 501.300 164.890 ;
        RECT 759.100 164.570 759.360 164.890 ;
        RECT 759.160 2.400 759.300 164.570 ;
        RECT 758.950 -4.800 759.510 2.400 ;
      LAYER via2 ;
        RECT 495.280 499.320 495.560 499.600 ;
        RECT 501.030 489.800 501.310 490.080 ;
      LAYER met3 ;
        RECT 495.255 499.620 495.585 499.625 ;
        RECT 495.230 499.610 495.610 499.620 ;
        RECT 494.800 499.310 495.610 499.610 ;
        RECT 495.230 499.300 495.610 499.310 ;
        RECT 495.255 499.295 495.585 499.300 ;
        RECT 495.230 490.090 495.610 490.100 ;
        RECT 501.005 490.090 501.335 490.105 ;
        RECT 495.230 489.790 501.335 490.090 ;
        RECT 495.230 489.780 495.610 489.790 ;
        RECT 501.005 489.775 501.335 489.790 ;
      LAYER via3 ;
        RECT 495.260 499.300 495.580 499.620 ;
        RECT 495.260 489.780 495.580 490.100 ;
      LAYER met4 ;
        RECT 495.255 499.295 495.585 499.625 ;
        RECT 495.270 490.105 495.570 499.295 ;
        RECT 495.255 489.775 495.585 490.105 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 596.000 499.500 596.320 499.760 ;
        RECT 596.090 499.080 596.230 499.500 ;
        RECT 595.770 498.880 596.230 499.080 ;
        RECT 595.770 498.820 596.090 498.880 ;
        RECT 595.770 493.580 596.090 493.640 ;
        RECT 597.150 493.580 597.470 493.640 ;
        RECT 595.770 493.440 597.470 493.580 ;
        RECT 595.770 493.380 596.090 493.440 ;
        RECT 597.150 493.380 597.470 493.440 ;
        RECT 597.150 162.760 597.470 162.820 ;
        RECT 2049.370 162.760 2049.690 162.820 ;
        RECT 597.150 162.620 2049.690 162.760 ;
        RECT 597.150 162.560 597.470 162.620 ;
        RECT 2049.370 162.560 2049.690 162.620 ;
      LAYER via ;
        RECT 596.030 499.500 596.290 499.760 ;
        RECT 595.800 498.820 596.060 499.080 ;
        RECT 595.800 493.380 596.060 493.640 ;
        RECT 597.180 493.380 597.440 493.640 ;
        RECT 597.180 162.560 597.440 162.820 ;
        RECT 2049.400 162.560 2049.660 162.820 ;
      LAYER met2 ;
        RECT 596.050 500.000 596.330 504.000 ;
        RECT 596.090 499.790 596.230 500.000 ;
        RECT 596.030 499.470 596.290 499.790 ;
        RECT 595.800 498.790 596.060 499.110 ;
        RECT 595.860 493.670 596.000 498.790 ;
        RECT 595.800 493.350 596.060 493.670 ;
        RECT 597.180 493.350 597.440 493.670 ;
        RECT 597.240 162.850 597.380 493.350 ;
        RECT 597.180 162.530 597.440 162.850 ;
        RECT 2049.400 162.530 2049.660 162.850 ;
        RECT 2049.460 82.870 2049.600 162.530 ;
        RECT 2049.460 82.730 2054.200 82.870 ;
        RECT 2054.060 2.400 2054.200 82.730 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 595.400 499.900 597.610 500.040 ;
        RECT 595.400 498.340 595.540 499.900 ;
        RECT 597.470 499.760 597.610 499.900 ;
        RECT 597.380 499.500 597.700 499.760 ;
        RECT 596.690 498.340 597.010 498.400 ;
        RECT 595.400 498.200 597.010 498.340 ;
        RECT 596.690 498.140 597.010 498.200 ;
        RECT 595.770 121.280 596.090 121.340 ;
        RECT 2070.070 121.280 2070.390 121.340 ;
        RECT 595.770 121.140 2070.390 121.280 ;
        RECT 595.770 121.080 596.090 121.140 ;
        RECT 2070.070 121.080 2070.390 121.140 ;
      LAYER via ;
        RECT 597.410 499.500 597.670 499.760 ;
        RECT 596.720 498.140 596.980 498.400 ;
        RECT 595.800 121.080 596.060 121.340 ;
        RECT 2070.100 121.080 2070.360 121.340 ;
      LAYER met2 ;
        RECT 597.430 500.000 597.710 504.000 ;
        RECT 597.470 499.790 597.610 500.000 ;
        RECT 597.410 499.470 597.670 499.790 ;
        RECT 596.720 498.110 596.980 498.430 ;
        RECT 596.780 473.010 596.920 498.110 ;
        RECT 595.860 472.870 596.920 473.010 ;
        RECT 595.860 121.370 596.000 472.870 ;
        RECT 595.800 121.050 596.060 121.370 ;
        RECT 2070.100 121.050 2070.360 121.370 ;
        RECT 2070.160 82.870 2070.300 121.050 ;
        RECT 2070.160 82.730 2071.680 82.870 ;
        RECT 2071.540 2.400 2071.680 82.730 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.810 500.000 599.090 504.000 ;
        RECT 598.850 498.680 598.990 500.000 ;
        RECT 598.620 498.540 598.990 498.680 ;
        RECT 598.620 497.605 598.760 498.540 ;
        RECT 598.550 497.235 598.830 497.605 ;
        RECT 2083.890 161.995 2084.170 162.365 ;
        RECT 2083.960 82.870 2084.100 161.995 ;
        RECT 2083.960 82.730 2087.320 82.870 ;
        RECT 2087.180 1.770 2087.320 82.730 ;
        RECT 2089.270 1.770 2089.830 2.400 ;
        RECT 2087.180 1.630 2089.830 1.770 ;
        RECT 2089.270 -4.800 2089.830 1.630 ;
      LAYER via2 ;
        RECT 598.550 497.280 598.830 497.560 ;
        RECT 2083.890 162.040 2084.170 162.320 ;
      LAYER met3 ;
        RECT 598.525 497.580 598.855 497.585 ;
        RECT 598.270 497.570 598.855 497.580 ;
        RECT 598.070 497.270 598.855 497.570 ;
        RECT 598.270 497.260 598.855 497.270 ;
        RECT 598.525 497.255 598.855 497.260 ;
        RECT 598.270 162.330 598.650 162.340 ;
        RECT 2083.865 162.330 2084.195 162.345 ;
        RECT 598.270 162.030 2084.195 162.330 ;
        RECT 598.270 162.020 598.650 162.030 ;
        RECT 2083.865 162.015 2084.195 162.030 ;
      LAYER via3 ;
        RECT 598.300 497.260 598.620 497.580 ;
        RECT 598.300 162.020 598.620 162.340 ;
      LAYER met4 ;
        RECT 598.295 497.255 598.625 497.585 ;
        RECT 598.310 162.345 598.610 497.255 ;
        RECT 598.295 162.015 598.625 162.345 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.140 499.500 600.460 499.760 ;
        RECT 600.230 498.400 600.370 499.500 ;
        RECT 600.230 498.200 600.690 498.400 ;
        RECT 600.370 498.140 600.690 498.200 ;
        RECT 600.830 471.820 601.150 471.880 ;
        RECT 602.210 471.820 602.530 471.880 ;
        RECT 600.830 471.680 602.530 471.820 ;
        RECT 600.830 471.620 601.150 471.680 ;
        RECT 602.210 471.620 602.530 471.680 ;
        RECT 602.210 162.420 602.530 162.480 ;
        RECT 2104.570 162.420 2104.890 162.480 ;
        RECT 602.210 162.280 2104.890 162.420 ;
        RECT 602.210 162.220 602.530 162.280 ;
        RECT 2104.570 162.220 2104.890 162.280 ;
      LAYER via ;
        RECT 600.170 499.500 600.430 499.760 ;
        RECT 600.400 498.140 600.660 498.400 ;
        RECT 600.860 471.620 601.120 471.880 ;
        RECT 602.240 471.620 602.500 471.880 ;
        RECT 602.240 162.220 602.500 162.480 ;
        RECT 2104.600 162.220 2104.860 162.480 ;
      LAYER met2 ;
        RECT 600.190 500.000 600.470 504.000 ;
        RECT 600.230 499.790 600.370 500.000 ;
        RECT 600.170 499.470 600.430 499.790 ;
        RECT 600.400 498.110 600.660 498.430 ;
        RECT 600.460 495.280 600.600 498.110 ;
        RECT 600.460 495.140 601.060 495.280 ;
        RECT 600.920 471.910 601.060 495.140 ;
        RECT 600.860 471.590 601.120 471.910 ;
        RECT 602.240 471.590 602.500 471.910 ;
        RECT 602.300 162.510 602.440 471.590 ;
        RECT 602.240 162.190 602.500 162.510 ;
        RECT 2104.600 162.190 2104.860 162.510 ;
        RECT 2104.660 1.770 2104.800 162.190 ;
        RECT 2106.750 1.770 2107.310 2.400 ;
        RECT 2104.660 1.630 2107.310 1.770 ;
        RECT 2106.750 -4.800 2107.310 1.630 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.370 65.860 600.690 65.920 ;
        RECT 2118.830 65.860 2119.150 65.920 ;
        RECT 600.370 65.720 2119.150 65.860 ;
        RECT 600.370 65.660 600.690 65.720 ;
        RECT 2118.830 65.660 2119.150 65.720 ;
        RECT 2118.830 16.900 2119.150 16.960 ;
        RECT 2124.810 16.900 2125.130 16.960 ;
        RECT 2118.830 16.760 2125.130 16.900 ;
        RECT 2118.830 16.700 2119.150 16.760 ;
        RECT 2124.810 16.700 2125.130 16.760 ;
      LAYER via ;
        RECT 600.400 65.660 600.660 65.920 ;
        RECT 2118.860 65.660 2119.120 65.920 ;
        RECT 2118.860 16.700 2119.120 16.960 ;
        RECT 2124.840 16.700 2125.100 16.960 ;
      LAYER met2 ;
        RECT 601.570 500.000 601.850 504.000 ;
        RECT 601.610 498.965 601.750 500.000 ;
        RECT 601.540 498.595 601.820 498.965 ;
        RECT 599.930 497.235 600.210 497.605 ;
        RECT 600.000 489.970 600.140 497.235 ;
        RECT 600.000 489.830 600.600 489.970 ;
        RECT 600.460 65.950 600.600 489.830 ;
        RECT 600.400 65.630 600.660 65.950 ;
        RECT 2118.860 65.630 2119.120 65.950 ;
        RECT 2118.920 16.990 2119.060 65.630 ;
        RECT 2118.860 16.670 2119.120 16.990 ;
        RECT 2124.840 16.670 2125.100 16.990 ;
        RECT 2124.900 2.400 2125.040 16.670 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
      LAYER via2 ;
        RECT 601.540 498.640 601.820 498.920 ;
        RECT 599.930 497.280 600.210 497.560 ;
      LAYER met3 ;
        RECT 601.515 498.615 601.845 498.945 ;
        RECT 599.905 497.570 600.235 497.585 ;
        RECT 601.530 497.570 601.830 498.615 ;
        RECT 599.905 497.270 601.830 497.570 ;
        RECT 599.905 497.255 600.235 497.270 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 602.900 499.500 603.220 499.760 ;
        RECT 602.990 498.400 603.130 499.500 ;
        RECT 602.670 498.200 603.130 498.400 ;
        RECT 602.670 498.140 602.990 498.200 ;
        RECT 601.750 472.840 602.070 472.900 ;
        RECT 602.670 472.840 602.990 472.900 ;
        RECT 601.750 472.700 602.990 472.840 ;
        RECT 601.750 472.640 602.070 472.700 ;
        RECT 602.670 472.640 602.990 472.700 ;
        RECT 601.750 114.820 602.070 114.880 ;
        RECT 2139.070 114.820 2139.390 114.880 ;
        RECT 601.750 114.680 2139.390 114.820 ;
        RECT 601.750 114.620 602.070 114.680 ;
        RECT 2139.070 114.620 2139.390 114.680 ;
      LAYER via ;
        RECT 602.930 499.500 603.190 499.760 ;
        RECT 602.700 498.140 602.960 498.400 ;
        RECT 601.780 472.640 602.040 472.900 ;
        RECT 602.700 472.640 602.960 472.900 ;
        RECT 601.780 114.620 602.040 114.880 ;
        RECT 2139.100 114.620 2139.360 114.880 ;
      LAYER met2 ;
        RECT 602.950 500.000 603.230 504.000 ;
        RECT 602.990 499.790 603.130 500.000 ;
        RECT 602.930 499.470 603.190 499.790 ;
        RECT 602.700 498.110 602.960 498.430 ;
        RECT 602.760 472.930 602.900 498.110 ;
        RECT 601.780 472.610 602.040 472.930 ;
        RECT 602.700 472.610 602.960 472.930 ;
        RECT 601.840 114.910 601.980 472.610 ;
        RECT 601.780 114.590 602.040 114.910 ;
        RECT 2139.100 114.590 2139.360 114.910 ;
        RECT 2139.160 82.870 2139.300 114.590 ;
        RECT 2139.160 82.730 2142.520 82.870 ;
        RECT 2142.380 2.400 2142.520 82.730 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 604.280 499.500 604.600 499.760 ;
        RECT 604.370 498.060 604.510 499.500 ;
        RECT 604.370 497.860 604.830 498.060 ;
        RECT 604.510 497.800 604.830 497.860 ;
        RECT 603.590 169.220 603.910 169.280 ;
        RECT 2159.770 169.220 2160.090 169.280 ;
        RECT 603.590 169.080 2160.090 169.220 ;
        RECT 603.590 169.020 603.910 169.080 ;
        RECT 2159.770 169.020 2160.090 169.080 ;
      LAYER via ;
        RECT 604.310 499.500 604.570 499.760 ;
        RECT 604.540 497.800 604.800 498.060 ;
        RECT 603.620 169.020 603.880 169.280 ;
        RECT 2159.800 169.020 2160.060 169.280 ;
      LAYER met2 ;
        RECT 604.330 500.000 604.610 504.000 ;
        RECT 604.370 499.790 604.510 500.000 ;
        RECT 604.310 499.470 604.570 499.790 ;
        RECT 604.540 497.770 604.800 498.090 ;
        RECT 604.600 496.130 604.740 497.770 ;
        RECT 604.140 495.990 604.740 496.130 ;
        RECT 604.140 420.970 604.280 495.990 ;
        RECT 603.680 420.830 604.280 420.970 ;
        RECT 603.680 169.310 603.820 420.830 ;
        RECT 603.620 168.990 603.880 169.310 ;
        RECT 2159.800 168.990 2160.060 169.310 ;
        RECT 2159.860 5.850 2160.000 168.990 ;
        RECT 2159.860 5.710 2160.460 5.850 ;
        RECT 2160.320 2.400 2160.460 5.710 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 605.660 499.500 605.980 499.760 ;
        RECT 605.750 499.360 605.890 499.500 ;
        RECT 605.520 499.220 605.890 499.360 ;
        RECT 605.520 498.680 605.660 499.220 ;
        RECT 606.350 498.680 606.670 498.740 ;
        RECT 605.520 498.540 606.670 498.680 ;
        RECT 606.350 498.480 606.670 498.540 ;
      LAYER via ;
        RECT 605.690 499.500 605.950 499.760 ;
        RECT 606.380 498.480 606.640 498.740 ;
      LAYER met2 ;
        RECT 605.710 500.000 605.990 504.000 ;
        RECT 605.750 499.790 605.890 500.000 ;
        RECT 605.690 499.470 605.950 499.790 ;
        RECT 606.380 498.450 606.640 498.770 ;
        RECT 606.440 491.485 606.580 498.450 ;
        RECT 606.370 491.115 606.650 491.485 ;
        RECT 2173.590 129.355 2173.870 129.725 ;
        RECT 2173.660 82.870 2173.800 129.355 ;
        RECT 2173.660 82.730 2175.640 82.870 ;
        RECT 2175.500 1.770 2175.640 82.730 ;
        RECT 2177.590 1.770 2178.150 2.400 ;
        RECT 2175.500 1.630 2178.150 1.770 ;
        RECT 2177.590 -4.800 2178.150 1.630 ;
      LAYER via2 ;
        RECT 606.370 491.160 606.650 491.440 ;
        RECT 2173.590 129.400 2173.870 129.680 ;
      LAYER met3 ;
        RECT 604.710 491.450 605.090 491.460 ;
        RECT 606.345 491.450 606.675 491.465 ;
        RECT 604.710 491.150 606.675 491.450 ;
        RECT 604.710 491.140 605.090 491.150 ;
        RECT 606.345 491.135 606.675 491.150 ;
        RECT 604.710 129.690 605.090 129.700 ;
        RECT 2173.565 129.690 2173.895 129.705 ;
        RECT 604.710 129.390 2173.895 129.690 ;
        RECT 604.710 129.380 605.090 129.390 ;
        RECT 2173.565 129.375 2173.895 129.390 ;
      LAYER via3 ;
        RECT 604.740 491.140 605.060 491.460 ;
        RECT 604.740 129.380 605.060 129.700 ;
      LAYER met4 ;
        RECT 604.735 491.135 605.065 491.465 ;
        RECT 604.750 129.705 605.050 491.135 ;
        RECT 604.735 129.375 605.065 129.705 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.040 498.820 607.360 499.080 ;
        RECT 607.130 498.060 607.270 498.820 ;
        RECT 606.810 497.860 607.270 498.060 ;
        RECT 606.810 497.800 607.130 497.860 ;
        RECT 607.270 472.840 607.590 472.900 ;
        RECT 609.570 472.840 609.890 472.900 ;
        RECT 607.270 472.700 609.890 472.840 ;
        RECT 607.270 472.640 607.590 472.700 ;
        RECT 609.570 472.640 609.890 472.700 ;
        RECT 609.570 136.580 609.890 136.640 ;
        RECT 2194.270 136.580 2194.590 136.640 ;
        RECT 609.570 136.440 2194.590 136.580 ;
        RECT 609.570 136.380 609.890 136.440 ;
        RECT 2194.270 136.380 2194.590 136.440 ;
      LAYER via ;
        RECT 607.070 498.820 607.330 499.080 ;
        RECT 606.840 497.800 607.100 498.060 ;
        RECT 607.300 472.640 607.560 472.900 ;
        RECT 609.600 472.640 609.860 472.900 ;
        RECT 609.600 136.380 609.860 136.640 ;
        RECT 2194.300 136.380 2194.560 136.640 ;
      LAYER met2 ;
        RECT 607.090 500.000 607.370 504.000 ;
        RECT 607.130 499.110 607.270 500.000 ;
        RECT 607.070 498.790 607.330 499.110 ;
        RECT 606.840 497.770 607.100 498.090 ;
        RECT 606.900 483.070 607.040 497.770 ;
        RECT 606.900 482.930 607.500 483.070 ;
        RECT 607.360 472.930 607.500 482.930 ;
        RECT 607.300 472.610 607.560 472.930 ;
        RECT 609.600 472.610 609.860 472.930 ;
        RECT 609.660 136.670 609.800 472.610 ;
        RECT 609.600 136.350 609.860 136.670 ;
        RECT 2194.300 136.350 2194.560 136.670 ;
        RECT 2194.360 82.870 2194.500 136.350 ;
        RECT 2194.360 82.730 2195.880 82.870 ;
        RECT 2195.740 2.400 2195.880 82.730 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 608.650 136.240 608.970 136.300 ;
        RECT 2208.070 136.240 2208.390 136.300 ;
        RECT 608.650 136.100 2208.390 136.240 ;
        RECT 608.650 136.040 608.970 136.100 ;
        RECT 2208.070 136.040 2208.390 136.100 ;
      LAYER via ;
        RECT 608.680 136.040 608.940 136.300 ;
        RECT 2208.100 136.040 2208.360 136.300 ;
      LAYER met2 ;
        RECT 608.470 500.000 608.750 504.000 ;
        RECT 608.510 498.680 608.650 500.000 ;
        RECT 608.510 498.540 608.880 498.680 ;
        RECT 608.740 136.330 608.880 498.540 ;
        RECT 608.680 136.010 608.940 136.330 ;
        RECT 2208.100 136.010 2208.360 136.330 ;
        RECT 2208.160 82.870 2208.300 136.010 ;
        RECT 2208.160 82.730 2213.360 82.870 ;
        RECT 2213.220 2.400 2213.360 82.730 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.640 499.160 496.960 499.420 ;
        RECT 496.730 498.680 496.870 499.160 ;
        RECT 496.500 498.540 496.870 498.680 ;
        RECT 496.500 496.300 496.640 498.540 ;
        RECT 497.330 496.300 497.650 496.360 ;
        RECT 496.500 496.160 497.650 496.300 ;
        RECT 497.330 496.100 497.650 496.160 ;
        RECT 497.330 473.520 497.650 473.580 ;
        RECT 497.330 473.380 500.320 473.520 ;
        RECT 497.330 473.320 497.650 473.380 ;
        RECT 499.630 472.160 499.950 472.220 ;
        RECT 500.180 472.160 500.320 473.380 ;
        RECT 499.630 472.020 500.320 472.160 ;
        RECT 499.630 471.960 499.950 472.020 ;
        RECT 499.630 130.460 499.950 130.520 ;
        RECT 772.870 130.460 773.190 130.520 ;
        RECT 499.630 130.320 773.190 130.460 ;
        RECT 499.630 130.260 499.950 130.320 ;
        RECT 772.870 130.260 773.190 130.320 ;
      LAYER via ;
        RECT 496.670 499.160 496.930 499.420 ;
        RECT 497.360 496.100 497.620 496.360 ;
        RECT 497.360 473.320 497.620 473.580 ;
        RECT 499.660 471.960 499.920 472.220 ;
        RECT 499.660 130.260 499.920 130.520 ;
        RECT 772.900 130.260 773.160 130.520 ;
      LAYER met2 ;
        RECT 496.690 500.000 496.970 504.000 ;
        RECT 496.730 499.450 496.870 500.000 ;
        RECT 496.670 499.130 496.930 499.450 ;
        RECT 497.360 496.070 497.620 496.390 ;
        RECT 497.420 473.610 497.560 496.070 ;
        RECT 497.360 473.290 497.620 473.610 ;
        RECT 499.660 471.930 499.920 472.250 ;
        RECT 499.720 130.550 499.860 471.930 ;
        RECT 499.660 130.230 499.920 130.550 ;
        RECT 772.900 130.230 773.160 130.550 ;
        RECT 772.960 82.870 773.100 130.230 ;
        RECT 772.960 82.730 777.240 82.870 ;
        RECT 777.100 2.400 777.240 82.730 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 609.800 499.160 610.120 499.420 ;
        RECT 609.890 498.340 610.030 499.160 ;
        RECT 609.200 498.200 610.030 498.340 ;
        RECT 609.200 497.720 609.340 498.200 ;
        RECT 609.110 497.460 609.430 497.720 ;
        RECT 609.110 135.900 609.430 135.960 ;
        RECT 2228.770 135.900 2229.090 135.960 ;
        RECT 609.110 135.760 2229.090 135.900 ;
        RECT 609.110 135.700 609.430 135.760 ;
        RECT 2228.770 135.700 2229.090 135.760 ;
      LAYER via ;
        RECT 609.830 499.160 610.090 499.420 ;
        RECT 609.140 497.460 609.400 497.720 ;
        RECT 609.140 135.700 609.400 135.960 ;
        RECT 2228.800 135.700 2229.060 135.960 ;
      LAYER met2 ;
        RECT 609.850 500.000 610.130 504.000 ;
        RECT 609.890 499.450 610.030 500.000 ;
        RECT 609.830 499.130 610.090 499.450 ;
        RECT 609.140 497.430 609.400 497.750 ;
        RECT 609.200 135.990 609.340 497.430 ;
        RECT 609.140 135.670 609.400 135.990 ;
        RECT 2228.800 135.670 2229.060 135.990 ;
        RECT 2228.860 1.770 2229.000 135.670 ;
        RECT 2230.950 1.770 2231.510 2.400 ;
        RECT 2228.860 1.630 2231.510 1.770 ;
        RECT 2230.950 -4.800 2231.510 1.630 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 611.180 499.160 611.500 499.420 ;
        RECT 611.270 498.340 611.410 499.160 ;
        RECT 611.870 498.340 612.190 498.400 ;
        RECT 611.270 498.200 612.190 498.340 ;
        RECT 611.870 498.140 612.190 498.200 ;
        RECT 607.270 472.160 607.590 472.220 ;
        RECT 611.870 472.160 612.190 472.220 ;
        RECT 607.270 472.020 612.190 472.160 ;
        RECT 607.270 471.960 607.590 472.020 ;
        RECT 611.870 471.960 612.190 472.020 ;
        RECT 607.270 94.080 607.590 94.140 ;
        RECT 2243.030 94.080 2243.350 94.140 ;
        RECT 607.270 93.940 2243.350 94.080 ;
        RECT 607.270 93.880 607.590 93.940 ;
        RECT 2243.030 93.880 2243.350 93.940 ;
        RECT 2243.030 16.900 2243.350 16.960 ;
        RECT 2249.010 16.900 2249.330 16.960 ;
        RECT 2243.030 16.760 2249.330 16.900 ;
        RECT 2243.030 16.700 2243.350 16.760 ;
        RECT 2249.010 16.700 2249.330 16.760 ;
      LAYER via ;
        RECT 611.210 499.160 611.470 499.420 ;
        RECT 611.900 498.140 612.160 498.400 ;
        RECT 607.300 471.960 607.560 472.220 ;
        RECT 611.900 471.960 612.160 472.220 ;
        RECT 607.300 93.880 607.560 94.140 ;
        RECT 2243.060 93.880 2243.320 94.140 ;
        RECT 2243.060 16.700 2243.320 16.960 ;
        RECT 2249.040 16.700 2249.300 16.960 ;
      LAYER met2 ;
        RECT 611.230 500.000 611.510 504.000 ;
        RECT 611.270 499.450 611.410 500.000 ;
        RECT 611.210 499.130 611.470 499.450 ;
        RECT 611.900 498.110 612.160 498.430 ;
        RECT 611.960 472.250 612.100 498.110 ;
        RECT 607.300 471.930 607.560 472.250 ;
        RECT 611.900 471.930 612.160 472.250 ;
        RECT 607.360 94.170 607.500 471.930 ;
        RECT 607.300 93.850 607.560 94.170 ;
        RECT 2243.060 93.850 2243.320 94.170 ;
        RECT 2243.120 16.990 2243.260 93.850 ;
        RECT 2243.060 16.670 2243.320 16.990 ;
        RECT 2249.040 16.670 2249.300 16.990 ;
        RECT 2249.100 2.400 2249.240 16.670 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 612.560 499.500 612.880 499.760 ;
        RECT 612.650 498.400 612.790 499.500 ;
        RECT 612.650 498.200 613.110 498.400 ;
        RECT 612.790 498.140 613.110 498.200 ;
      LAYER via ;
        RECT 612.590 499.500 612.850 499.760 ;
        RECT 612.820 498.140 613.080 498.400 ;
      LAYER met2 ;
        RECT 612.610 500.000 612.890 504.000 ;
        RECT 612.650 499.790 612.790 500.000 ;
        RECT 612.590 499.470 612.850 499.790 ;
        RECT 612.820 498.110 613.080 498.430 ;
        RECT 612.880 484.685 613.020 498.110 ;
        RECT 612.810 484.315 613.090 484.685 ;
        RECT 2263.290 168.795 2263.570 169.165 ;
        RECT 2263.360 82.870 2263.500 168.795 ;
        RECT 2263.360 82.730 2266.720 82.870 ;
        RECT 2266.580 2.400 2266.720 82.730 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
      LAYER via2 ;
        RECT 612.810 484.360 613.090 484.640 ;
        RECT 2263.290 168.840 2263.570 169.120 ;
      LAYER met3 ;
        RECT 611.150 484.650 611.530 484.660 ;
        RECT 612.785 484.650 613.115 484.665 ;
        RECT 611.150 484.350 613.115 484.650 ;
        RECT 611.150 484.340 611.530 484.350 ;
        RECT 612.785 484.335 613.115 484.350 ;
        RECT 611.150 169.130 611.530 169.140 ;
        RECT 2263.265 169.130 2263.595 169.145 ;
        RECT 611.150 168.830 2263.595 169.130 ;
        RECT 611.150 168.820 611.530 168.830 ;
        RECT 2263.265 168.815 2263.595 168.830 ;
      LAYER via3 ;
        RECT 611.180 484.340 611.500 484.660 ;
        RECT 611.180 168.820 611.500 169.140 ;
      LAYER met4 ;
        RECT 611.175 484.335 611.505 484.665 ;
        RECT 611.190 169.145 611.490 484.335 ;
        RECT 611.175 168.815 611.505 169.145 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 613.940 499.360 614.260 499.420 ;
        RECT 613.940 499.220 615.320 499.360 ;
        RECT 613.940 499.160 614.260 499.220 ;
        RECT 615.180 498.740 615.320 499.220 ;
        RECT 615.090 498.480 615.410 498.740 ;
        RECT 615.550 128.420 615.870 128.480 ;
        RECT 2284.430 128.420 2284.750 128.480 ;
        RECT 615.550 128.280 2284.750 128.420 ;
        RECT 615.550 128.220 615.870 128.280 ;
        RECT 2284.430 128.220 2284.750 128.280 ;
      LAYER via ;
        RECT 613.970 499.160 614.230 499.420 ;
        RECT 615.120 498.480 615.380 498.740 ;
        RECT 615.580 128.220 615.840 128.480 ;
        RECT 2284.460 128.220 2284.720 128.480 ;
      LAYER met2 ;
        RECT 613.990 500.000 614.270 504.000 ;
        RECT 614.030 499.450 614.170 500.000 ;
        RECT 613.970 499.130 614.230 499.450 ;
        RECT 615.120 498.450 615.380 498.770 ;
        RECT 615.180 479.130 615.320 498.450 ;
        RECT 615.180 478.990 615.780 479.130 ;
        RECT 615.640 128.510 615.780 478.990 ;
        RECT 615.580 128.190 615.840 128.510 ;
        RECT 2284.460 128.190 2284.720 128.510 ;
        RECT 2284.520 2.400 2284.660 128.190 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 615.550 479.640 615.870 479.700 ;
        RECT 616.930 479.640 617.250 479.700 ;
        RECT 615.550 479.500 617.250 479.640 ;
        RECT 615.550 479.440 615.870 479.500 ;
        RECT 616.930 479.440 617.250 479.500 ;
        RECT 616.930 168.880 617.250 168.940 ;
        RECT 2297.770 168.880 2298.090 168.940 ;
        RECT 616.930 168.740 2298.090 168.880 ;
        RECT 616.930 168.680 617.250 168.740 ;
        RECT 2297.770 168.680 2298.090 168.740 ;
      LAYER via ;
        RECT 615.580 479.440 615.840 479.700 ;
        RECT 616.960 479.440 617.220 479.700 ;
        RECT 616.960 168.680 617.220 168.940 ;
        RECT 2297.800 168.680 2298.060 168.940 ;
      LAYER met2 ;
        RECT 615.370 500.000 615.650 504.000 ;
        RECT 615.410 499.360 615.550 500.000 ;
        RECT 615.410 499.220 615.780 499.360 ;
        RECT 615.640 479.730 615.780 499.220 ;
        RECT 615.580 479.410 615.840 479.730 ;
        RECT 616.960 479.410 617.220 479.730 ;
        RECT 617.020 168.970 617.160 479.410 ;
        RECT 616.960 168.650 617.220 168.970 ;
        RECT 2297.800 168.650 2298.060 168.970 ;
        RECT 2297.860 82.870 2298.000 168.650 ;
        RECT 2297.860 82.730 2299.840 82.870 ;
        RECT 2299.700 1.770 2299.840 82.730 ;
        RECT 2301.790 1.770 2302.350 2.400 ;
        RECT 2299.700 1.630 2302.350 1.770 ;
        RECT 2301.790 -4.800 2302.350 1.630 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 616.700 499.160 617.020 499.420 ;
        RECT 616.010 498.340 616.330 498.400 ;
        RECT 616.790 498.340 616.930 499.160 ;
        RECT 616.010 498.200 616.930 498.340 ;
        RECT 616.010 498.140 616.330 498.200 ;
        RECT 616.010 135.560 616.330 135.620 ;
        RECT 2318.470 135.560 2318.790 135.620 ;
        RECT 616.010 135.420 2318.790 135.560 ;
        RECT 616.010 135.360 616.330 135.420 ;
        RECT 2318.470 135.360 2318.790 135.420 ;
      LAYER via ;
        RECT 616.730 499.160 616.990 499.420 ;
        RECT 616.040 498.140 616.300 498.400 ;
        RECT 616.040 135.360 616.300 135.620 ;
        RECT 2318.500 135.360 2318.760 135.620 ;
      LAYER met2 ;
        RECT 616.750 500.000 617.030 504.000 ;
        RECT 616.790 499.450 616.930 500.000 ;
        RECT 616.730 499.130 616.990 499.450 ;
        RECT 616.040 498.110 616.300 498.430 ;
        RECT 616.100 135.650 616.240 498.110 ;
        RECT 616.040 135.330 616.300 135.650 ;
        RECT 2318.500 135.330 2318.760 135.650 ;
        RECT 2318.560 82.870 2318.700 135.330 ;
        RECT 2318.560 82.730 2320.080 82.870 ;
        RECT 2319.940 2.400 2320.080 82.730 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 616.470 472.840 616.790 472.900 ;
        RECT 618.310 472.840 618.630 472.900 ;
        RECT 616.470 472.700 618.630 472.840 ;
        RECT 616.470 472.640 616.790 472.700 ;
        RECT 618.310 472.640 618.630 472.700 ;
        RECT 616.470 149.500 616.790 149.560 ;
        RECT 2332.270 149.500 2332.590 149.560 ;
        RECT 616.470 149.360 2332.590 149.500 ;
        RECT 616.470 149.300 616.790 149.360 ;
        RECT 2332.270 149.300 2332.590 149.360 ;
      LAYER via ;
        RECT 616.500 472.640 616.760 472.900 ;
        RECT 618.340 472.640 618.600 472.900 ;
        RECT 616.500 149.300 616.760 149.560 ;
        RECT 2332.300 149.300 2332.560 149.560 ;
      LAYER met2 ;
        RECT 618.130 500.000 618.410 504.000 ;
        RECT 618.170 498.680 618.310 500.000 ;
        RECT 618.170 498.540 618.540 498.680 ;
        RECT 618.400 472.930 618.540 498.540 ;
        RECT 616.500 472.610 616.760 472.930 ;
        RECT 618.340 472.610 618.600 472.930 ;
        RECT 616.560 149.590 616.700 472.610 ;
        RECT 616.500 149.270 616.760 149.590 ;
        RECT 2332.300 149.270 2332.560 149.590 ;
        RECT 2332.360 82.870 2332.500 149.270 ;
        RECT 2332.360 82.730 2337.560 82.870 ;
        RECT 2337.420 2.400 2337.560 82.730 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 614.630 473.180 614.950 473.240 ;
        RECT 619.690 473.180 620.010 473.240 ;
        RECT 614.630 473.040 620.010 473.180 ;
        RECT 614.630 472.980 614.950 473.040 ;
        RECT 619.690 472.980 620.010 473.040 ;
        RECT 614.630 93.740 614.950 93.800 ;
        RECT 2352.970 93.740 2353.290 93.800 ;
        RECT 614.630 93.600 2353.290 93.740 ;
        RECT 614.630 93.540 614.950 93.600 ;
        RECT 2352.970 93.540 2353.290 93.600 ;
      LAYER via ;
        RECT 614.660 472.980 614.920 473.240 ;
        RECT 619.720 472.980 619.980 473.240 ;
        RECT 614.660 93.540 614.920 93.800 ;
        RECT 2353.000 93.540 2353.260 93.800 ;
      LAYER met2 ;
        RECT 619.510 500.000 619.790 504.000 ;
        RECT 619.550 498.340 619.690 500.000 ;
        RECT 619.550 498.200 619.920 498.340 ;
        RECT 619.780 473.270 619.920 498.200 ;
        RECT 614.660 472.950 614.920 473.270 ;
        RECT 619.720 472.950 619.980 473.270 ;
        RECT 614.720 93.830 614.860 472.950 ;
        RECT 614.660 93.510 614.920 93.830 ;
        RECT 2353.000 93.510 2353.260 93.830 ;
        RECT 2353.060 1.770 2353.200 93.510 ;
        RECT 2355.150 1.770 2355.710 2.400 ;
        RECT 2353.060 1.630 2355.710 1.770 ;
        RECT 2355.150 -4.800 2355.710 1.630 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 620.840 499.500 621.160 499.760 ;
        RECT 620.930 499.080 621.070 499.500 ;
        RECT 620.610 498.880 621.070 499.080 ;
        RECT 620.610 498.820 620.930 498.880 ;
        RECT 620.610 491.540 620.930 491.600 ;
        RECT 623.830 491.540 624.150 491.600 ;
        RECT 620.610 491.400 624.150 491.540 ;
        RECT 620.610 491.340 620.930 491.400 ;
        RECT 623.830 491.340 624.150 491.400 ;
        RECT 623.830 135.220 624.150 135.280 ;
        RECT 2366.770 135.220 2367.090 135.280 ;
        RECT 623.830 135.080 2367.090 135.220 ;
        RECT 623.830 135.020 624.150 135.080 ;
        RECT 2366.770 135.020 2367.090 135.080 ;
        RECT 2366.770 16.900 2367.090 16.960 ;
        RECT 2370.910 16.900 2371.230 16.960 ;
        RECT 2366.770 16.760 2371.230 16.900 ;
        RECT 2366.770 16.700 2367.090 16.760 ;
        RECT 2370.910 16.700 2371.230 16.760 ;
      LAYER via ;
        RECT 620.870 499.500 621.130 499.760 ;
        RECT 620.640 498.820 620.900 499.080 ;
        RECT 620.640 491.340 620.900 491.600 ;
        RECT 623.860 491.340 624.120 491.600 ;
        RECT 623.860 135.020 624.120 135.280 ;
        RECT 2366.800 135.020 2367.060 135.280 ;
        RECT 2366.800 16.700 2367.060 16.960 ;
        RECT 2370.940 16.700 2371.200 16.960 ;
      LAYER met2 ;
        RECT 620.890 500.000 621.170 504.000 ;
        RECT 620.930 499.790 621.070 500.000 ;
        RECT 620.870 499.470 621.130 499.790 ;
        RECT 620.640 498.790 620.900 499.110 ;
        RECT 620.700 491.630 620.840 498.790 ;
        RECT 620.640 491.310 620.900 491.630 ;
        RECT 623.860 491.310 624.120 491.630 ;
        RECT 623.920 135.310 624.060 491.310 ;
        RECT 623.860 134.990 624.120 135.310 ;
        RECT 2366.800 134.990 2367.060 135.310 ;
        RECT 2366.860 16.990 2367.000 134.990 ;
        RECT 2366.800 16.670 2367.060 16.990 ;
        RECT 2370.940 16.670 2371.200 16.990 ;
        RECT 2371.000 1.770 2371.140 16.670 ;
        RECT 2372.630 1.770 2373.190 2.400 ;
        RECT 2371.000 1.630 2373.190 1.770 ;
        RECT 2372.630 -4.800 2373.190 1.630 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.310 499.900 624.980 500.040 ;
        RECT 622.310 499.760 622.450 499.900 ;
        RECT 622.220 499.500 622.540 499.760 ;
        RECT 624.840 497.720 624.980 499.900 ;
        RECT 624.750 497.460 625.070 497.720 ;
        RECT 624.290 134.880 624.610 134.940 ;
        RECT 2387.470 134.880 2387.790 134.940 ;
        RECT 624.290 134.740 2387.790 134.880 ;
        RECT 624.290 134.680 624.610 134.740 ;
        RECT 2387.470 134.680 2387.790 134.740 ;
      LAYER via ;
        RECT 622.250 499.500 622.510 499.760 ;
        RECT 624.780 497.460 625.040 497.720 ;
        RECT 624.320 134.680 624.580 134.940 ;
        RECT 2387.500 134.680 2387.760 134.940 ;
      LAYER met2 ;
        RECT 622.270 500.000 622.550 504.000 ;
        RECT 622.310 499.790 622.450 500.000 ;
        RECT 622.250 499.470 622.510 499.790 ;
        RECT 624.780 497.430 625.040 497.750 ;
        RECT 624.840 473.010 624.980 497.430 ;
        RECT 624.380 472.870 624.980 473.010 ;
        RECT 624.380 134.970 624.520 472.870 ;
        RECT 624.320 134.650 624.580 134.970 ;
        RECT 2387.500 134.650 2387.760 134.970 ;
        RECT 2387.560 82.870 2387.700 134.650 ;
        RECT 2387.560 82.730 2390.920 82.870 ;
        RECT 2390.780 2.400 2390.920 82.730 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 498.020 499.500 498.340 499.760 ;
        RECT 498.110 499.080 498.250 499.500 ;
        RECT 498.020 498.820 498.340 499.080 ;
        RECT 498.250 95.780 498.570 95.840 ;
        RECT 793.570 95.780 793.890 95.840 ;
        RECT 498.250 95.640 793.890 95.780 ;
        RECT 498.250 95.580 498.570 95.640 ;
        RECT 793.570 95.580 793.890 95.640 ;
      LAYER via ;
        RECT 498.050 499.500 498.310 499.760 ;
        RECT 498.050 498.820 498.310 499.080 ;
        RECT 498.280 95.580 498.540 95.840 ;
        RECT 793.600 95.580 793.860 95.840 ;
      LAYER met2 ;
        RECT 498.070 500.000 498.350 504.000 ;
        RECT 498.110 499.790 498.250 500.000 ;
        RECT 498.050 499.470 498.310 499.790 ;
        RECT 498.050 498.790 498.310 499.110 ;
        RECT 498.110 498.340 498.250 498.790 ;
        RECT 498.110 498.200 498.480 498.340 ;
        RECT 498.340 95.870 498.480 498.200 ;
        RECT 498.280 95.550 498.540 95.870 ;
        RECT 793.600 95.550 793.860 95.870 ;
        RECT 793.660 82.870 793.800 95.550 ;
        RECT 793.660 82.730 794.720 82.870 ;
        RECT 794.580 2.400 794.720 82.730 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.070 498.340 483.390 498.400 ;
        RECT 485.830 498.340 486.150 498.400 ;
        RECT 483.070 498.200 486.150 498.340 ;
        RECT 483.070 498.140 483.390 498.200 ;
        RECT 485.830 498.140 486.150 498.200 ;
        RECT 541.490 19.620 541.810 19.680 ;
        RECT 640.850 19.620 641.170 19.680 ;
        RECT 541.490 19.480 641.170 19.620 ;
        RECT 541.490 19.420 541.810 19.480 ;
        RECT 640.850 19.420 641.170 19.480 ;
        RECT 483.530 18.260 483.850 18.320 ;
        RECT 541.490 18.260 541.810 18.320 ;
        RECT 483.530 18.120 541.810 18.260 ;
        RECT 483.530 18.060 483.850 18.120 ;
        RECT 541.490 18.060 541.810 18.120 ;
      LAYER via ;
        RECT 483.100 498.140 483.360 498.400 ;
        RECT 485.860 498.140 486.120 498.400 ;
        RECT 541.520 19.420 541.780 19.680 ;
        RECT 640.880 19.420 641.140 19.680 ;
        RECT 483.560 18.060 483.820 18.320 ;
        RECT 541.520 18.060 541.780 18.320 ;
      LAYER met2 ;
        RECT 486.110 500.000 486.390 504.000 ;
        RECT 486.150 499.020 486.290 500.000 ;
        RECT 485.920 498.880 486.290 499.020 ;
        RECT 485.920 498.430 486.060 498.880 ;
        RECT 483.100 498.110 483.360 498.430 ;
        RECT 485.860 498.110 486.120 498.430 ;
        RECT 483.160 448.570 483.300 498.110 ;
        RECT 483.160 448.430 483.760 448.570 ;
        RECT 483.620 18.350 483.760 448.430 ;
        RECT 541.520 19.390 541.780 19.710 ;
        RECT 640.880 19.390 641.140 19.710 ;
        RECT 541.580 18.350 541.720 19.390 ;
        RECT 483.560 18.030 483.820 18.350 ;
        RECT 541.520 18.030 541.780 18.350 ;
        RECT 640.940 2.400 641.080 19.390 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.910 79.800 623.230 79.860 ;
        RECT 2411.850 79.800 2412.170 79.860 ;
        RECT 622.910 79.660 2412.170 79.800 ;
        RECT 622.910 79.600 623.230 79.660 ;
        RECT 2411.850 79.600 2412.170 79.660 ;
      LAYER via ;
        RECT 622.940 79.600 623.200 79.860 ;
        RECT 2411.880 79.600 2412.140 79.860 ;
      LAYER met2 ;
        RECT 624.110 500.000 624.390 504.000 ;
        RECT 624.150 499.020 624.290 500.000 ;
        RECT 623.000 498.880 624.290 499.020 ;
        RECT 623.000 79.890 623.140 498.880 ;
        RECT 622.940 79.570 623.200 79.890 ;
        RECT 2411.880 79.570 2412.140 79.890 ;
        RECT 2411.940 1.770 2412.080 79.570 ;
        RECT 2414.030 1.770 2414.590 2.400 ;
        RECT 2411.940 1.630 2414.590 1.770 ;
        RECT 2414.030 -4.800 2414.590 1.630 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 625.440 499.020 625.760 499.080 ;
        RECT 625.300 498.820 625.760 499.020 ;
        RECT 625.300 497.720 625.440 498.820 ;
        RECT 625.210 497.460 625.530 497.720 ;
        RECT 623.370 472.160 623.690 472.220 ;
        RECT 625.210 472.160 625.530 472.220 ;
        RECT 623.370 472.020 625.530 472.160 ;
        RECT 623.370 471.960 623.690 472.020 ;
        RECT 625.210 471.960 625.530 472.020 ;
        RECT 623.370 93.400 623.690 93.460 ;
        RECT 2428.870 93.400 2429.190 93.460 ;
        RECT 623.370 93.260 2429.190 93.400 ;
        RECT 623.370 93.200 623.690 93.260 ;
        RECT 2428.870 93.200 2429.190 93.260 ;
      LAYER via ;
        RECT 625.470 498.820 625.730 499.080 ;
        RECT 625.240 497.460 625.500 497.720 ;
        RECT 623.400 471.960 623.660 472.220 ;
        RECT 625.240 471.960 625.500 472.220 ;
        RECT 623.400 93.200 623.660 93.460 ;
        RECT 2428.900 93.200 2429.160 93.460 ;
      LAYER met2 ;
        RECT 625.490 500.000 625.770 504.000 ;
        RECT 625.530 499.110 625.670 500.000 ;
        RECT 625.470 498.790 625.730 499.110 ;
        RECT 625.240 497.430 625.500 497.750 ;
        RECT 625.300 472.250 625.440 497.430 ;
        RECT 623.400 471.930 623.660 472.250 ;
        RECT 625.240 471.930 625.500 472.250 ;
        RECT 623.460 93.490 623.600 471.930 ;
        RECT 623.400 93.170 623.660 93.490 ;
        RECT 2428.900 93.170 2429.160 93.490 ;
        RECT 2428.960 82.870 2429.100 93.170 ;
        RECT 2428.960 82.730 2432.320 82.870 ;
        RECT 2432.180 2.400 2432.320 82.730 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 626.820 499.160 627.140 499.420 ;
        RECT 625.670 496.980 625.990 497.040 ;
        RECT 626.910 496.980 627.050 499.160 ;
        RECT 625.670 496.840 627.050 496.980 ;
        RECT 625.670 496.780 625.990 496.840 ;
      LAYER via ;
        RECT 626.850 499.160 627.110 499.420 ;
        RECT 625.700 496.780 625.960 497.040 ;
      LAYER met2 ;
        RECT 626.870 500.000 627.150 504.000 ;
        RECT 626.910 499.450 627.050 500.000 ;
        RECT 626.850 499.130 627.110 499.450 ;
        RECT 625.700 496.750 625.960 497.070 ;
        RECT 625.760 483.325 625.900 496.750 ;
        RECT 625.690 482.955 625.970 483.325 ;
        RECT 2449.590 134.795 2449.870 135.165 ;
        RECT 2449.660 2.400 2449.800 134.795 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
      LAYER via2 ;
        RECT 625.690 483.000 625.970 483.280 ;
        RECT 2449.590 134.840 2449.870 135.120 ;
      LAYER met3 ;
        RECT 624.030 483.290 624.410 483.300 ;
        RECT 625.665 483.290 625.995 483.305 ;
        RECT 624.030 482.990 625.995 483.290 ;
        RECT 624.030 482.980 624.410 482.990 ;
        RECT 625.665 482.975 625.995 482.990 ;
        RECT 624.030 135.130 624.410 135.140 ;
        RECT 2449.565 135.130 2449.895 135.145 ;
        RECT 624.030 134.830 2449.895 135.130 ;
        RECT 624.030 134.820 624.410 134.830 ;
        RECT 2449.565 134.815 2449.895 134.830 ;
      LAYER via3 ;
        RECT 624.060 482.980 624.380 483.300 ;
        RECT 624.060 134.820 624.380 135.140 ;
      LAYER met4 ;
        RECT 624.055 482.975 624.385 483.305 ;
        RECT 624.070 135.145 624.370 482.975 ;
        RECT 624.055 134.815 624.385 135.145 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 630.730 93.060 631.050 93.120 ;
        RECT 2463.370 93.060 2463.690 93.120 ;
        RECT 630.730 92.920 2463.690 93.060 ;
        RECT 630.730 92.860 631.050 92.920 ;
        RECT 2463.370 92.860 2463.690 92.920 ;
      LAYER via ;
        RECT 630.760 92.860 631.020 93.120 ;
        RECT 2463.400 92.860 2463.660 93.120 ;
      LAYER met2 ;
        RECT 628.250 500.000 628.530 504.000 ;
        RECT 628.290 499.645 628.430 500.000 ;
        RECT 628.220 499.275 628.500 499.645 ;
        RECT 630.750 497.915 631.030 498.285 ;
        RECT 630.820 93.150 630.960 497.915 ;
        RECT 630.760 92.830 631.020 93.150 ;
        RECT 2463.400 92.830 2463.660 93.150 ;
        RECT 2463.460 82.870 2463.600 92.830 ;
        RECT 2463.460 82.730 2465.440 82.870 ;
        RECT 2465.300 1.770 2465.440 82.730 ;
        RECT 2467.390 1.770 2467.950 2.400 ;
        RECT 2465.300 1.630 2467.950 1.770 ;
        RECT 2467.390 -4.800 2467.950 1.630 ;
      LAYER via2 ;
        RECT 628.220 499.320 628.500 499.600 ;
        RECT 630.750 497.960 631.030 498.240 ;
      LAYER met3 ;
        RECT 628.195 499.610 628.525 499.625 ;
        RECT 628.195 499.310 630.810 499.610 ;
        RECT 628.195 499.295 628.525 499.310 ;
        RECT 630.510 498.265 630.810 499.310 ;
        RECT 630.510 497.950 631.055 498.265 ;
        RECT 630.725 497.935 631.055 497.950 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 629.580 499.160 629.900 499.420 ;
        RECT 629.670 498.000 629.810 499.160 ;
        RECT 631.190 498.000 631.510 498.060 ;
        RECT 629.670 497.860 631.510 498.000 ;
        RECT 631.190 497.800 631.510 497.860 ;
        RECT 631.190 142.700 631.510 142.760 ;
        RECT 2484.070 142.700 2484.390 142.760 ;
        RECT 631.190 142.560 2484.390 142.700 ;
        RECT 631.190 142.500 631.510 142.560 ;
        RECT 2484.070 142.500 2484.390 142.560 ;
      LAYER via ;
        RECT 629.610 499.160 629.870 499.420 ;
        RECT 631.220 497.800 631.480 498.060 ;
        RECT 631.220 142.500 631.480 142.760 ;
        RECT 2484.100 142.500 2484.360 142.760 ;
      LAYER met2 ;
        RECT 629.630 500.000 629.910 504.000 ;
        RECT 629.670 499.450 629.810 500.000 ;
        RECT 629.610 499.130 629.870 499.450 ;
        RECT 631.220 497.770 631.480 498.090 ;
        RECT 631.280 142.790 631.420 497.770 ;
        RECT 631.220 142.470 631.480 142.790 ;
        RECT 2484.100 142.470 2484.360 142.790 ;
        RECT 2484.160 82.870 2484.300 142.470 ;
        RECT 2484.160 82.730 2485.680 82.870 ;
        RECT 2485.540 2.400 2485.680 82.730 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 631.650 142.360 631.970 142.420 ;
        RECT 2497.870 142.360 2498.190 142.420 ;
        RECT 631.650 142.220 2498.190 142.360 ;
        RECT 631.650 142.160 631.970 142.220 ;
        RECT 2497.870 142.160 2498.190 142.220 ;
      LAYER via ;
        RECT 631.680 142.160 631.940 142.420 ;
        RECT 2497.900 142.160 2498.160 142.420 ;
      LAYER met2 ;
        RECT 631.010 500.000 631.290 504.000 ;
        RECT 631.050 498.680 631.190 500.000 ;
        RECT 631.050 498.540 631.880 498.680 ;
        RECT 631.740 142.450 631.880 498.540 ;
        RECT 631.680 142.130 631.940 142.450 ;
        RECT 2497.900 142.130 2498.160 142.450 ;
        RECT 2497.960 82.870 2498.100 142.130 ;
        RECT 2497.960 82.730 2503.160 82.870 ;
        RECT 2503.020 2.400 2503.160 82.730 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.390 500.000 632.670 504.000 ;
        RECT 632.430 498.680 632.570 500.000 ;
        RECT 632.200 498.540 632.570 498.680 ;
        RECT 632.200 483.325 632.340 498.540 ;
        RECT 632.130 482.955 632.410 483.325 ;
        RECT 2518.590 142.275 2518.870 142.645 ;
        RECT 2518.660 1.770 2518.800 142.275 ;
        RECT 2520.750 1.770 2521.310 2.400 ;
        RECT 2518.660 1.630 2521.310 1.770 ;
        RECT 2520.750 -4.800 2521.310 1.630 ;
      LAYER via2 ;
        RECT 632.130 483.000 632.410 483.280 ;
        RECT 2518.590 142.320 2518.870 142.600 ;
      LAYER met3 ;
        RECT 631.390 483.290 631.770 483.300 ;
        RECT 632.105 483.290 632.435 483.305 ;
        RECT 631.390 482.990 632.435 483.290 ;
        RECT 631.390 482.980 631.770 482.990 ;
        RECT 632.105 482.975 632.435 482.990 ;
        RECT 631.390 142.610 631.770 142.620 ;
        RECT 2518.565 142.610 2518.895 142.625 ;
        RECT 631.390 142.310 2518.895 142.610 ;
        RECT 631.390 142.300 631.770 142.310 ;
        RECT 2518.565 142.295 2518.895 142.310 ;
      LAYER via3 ;
        RECT 631.420 482.980 631.740 483.300 ;
        RECT 631.420 142.300 631.740 142.620 ;
      LAYER met4 ;
        RECT 631.415 482.975 631.745 483.305 ;
        RECT 631.430 142.625 631.730 482.975 ;
        RECT 631.415 142.295 631.745 142.625 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 633.720 499.160 634.040 499.420 ;
        RECT 632.570 497.660 632.890 497.720 ;
        RECT 633.810 497.660 633.950 499.160 ;
        RECT 632.570 497.520 633.950 497.660 ;
        RECT 632.570 497.460 632.890 497.520 ;
        RECT 2532.370 17.580 2532.690 17.640 ;
        RECT 2536.510 17.580 2536.830 17.640 ;
        RECT 2532.370 17.440 2536.830 17.580 ;
        RECT 2532.370 17.380 2532.690 17.440 ;
        RECT 2536.510 17.380 2536.830 17.440 ;
      LAYER via ;
        RECT 633.750 499.160 634.010 499.420 ;
        RECT 632.600 497.460 632.860 497.720 ;
        RECT 2532.400 17.380 2532.660 17.640 ;
        RECT 2536.540 17.380 2536.800 17.640 ;
      LAYER met2 ;
        RECT 633.770 500.000 634.050 504.000 ;
        RECT 633.810 499.450 633.950 500.000 ;
        RECT 633.750 499.130 634.010 499.450 ;
        RECT 632.600 497.430 632.860 497.750 ;
        RECT 632.660 491.485 632.800 497.430 ;
        RECT 632.590 491.115 632.870 491.485 ;
        RECT 2532.390 92.635 2532.670 93.005 ;
        RECT 2532.460 17.670 2532.600 92.635 ;
        RECT 2532.400 17.350 2532.660 17.670 ;
        RECT 2536.540 17.350 2536.800 17.670 ;
        RECT 2536.600 1.770 2536.740 17.350 ;
        RECT 2538.230 1.770 2538.790 2.400 ;
        RECT 2536.600 1.630 2538.790 1.770 ;
        RECT 2538.230 -4.800 2538.790 1.630 ;
      LAYER via2 ;
        RECT 632.590 491.160 632.870 491.440 ;
        RECT 2532.390 92.680 2532.670 92.960 ;
      LAYER met3 ;
        RECT 632.565 491.460 632.895 491.465 ;
        RECT 632.310 491.450 632.895 491.460 ;
        RECT 632.110 491.150 632.895 491.450 ;
        RECT 632.310 491.140 632.895 491.150 ;
        RECT 632.565 491.135 632.895 491.140 ;
        RECT 632.310 92.970 632.690 92.980 ;
        RECT 2532.365 92.970 2532.695 92.985 ;
        RECT 632.310 92.670 2532.695 92.970 ;
        RECT 632.310 92.660 632.690 92.670 ;
        RECT 2532.365 92.655 2532.695 92.670 ;
      LAYER via3 ;
        RECT 632.340 491.140 632.660 491.460 ;
        RECT 632.340 92.660 632.660 92.980 ;
      LAYER met4 ;
        RECT 632.335 491.135 632.665 491.465 ;
        RECT 632.350 92.985 632.650 491.135 ;
        RECT 632.335 92.655 632.665 92.985 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.870 471.820 635.190 471.880 ;
        RECT 637.170 471.820 637.490 471.880 ;
        RECT 634.870 471.680 637.490 471.820 ;
        RECT 634.870 471.620 635.190 471.680 ;
        RECT 637.170 471.620 637.490 471.680 ;
        RECT 637.170 134.540 637.490 134.600 ;
        RECT 2553.070 134.540 2553.390 134.600 ;
        RECT 637.170 134.400 2553.390 134.540 ;
        RECT 637.170 134.340 637.490 134.400 ;
        RECT 2553.070 134.340 2553.390 134.400 ;
      LAYER via ;
        RECT 634.900 471.620 635.160 471.880 ;
        RECT 637.200 471.620 637.460 471.880 ;
        RECT 637.200 134.340 637.460 134.600 ;
        RECT 2553.100 134.340 2553.360 134.600 ;
      LAYER met2 ;
        RECT 635.150 500.000 635.430 504.000 ;
        RECT 635.190 499.530 635.330 500.000 ;
        RECT 635.190 499.390 635.560 499.530 ;
        RECT 635.420 498.680 635.560 499.390 ;
        RECT 634.960 498.540 635.560 498.680 ;
        RECT 634.960 471.910 635.100 498.540 ;
        RECT 634.900 471.590 635.160 471.910 ;
        RECT 637.200 471.590 637.460 471.910 ;
        RECT 637.260 134.630 637.400 471.590 ;
        RECT 637.200 134.310 637.460 134.630 ;
        RECT 2553.100 134.310 2553.360 134.630 ;
        RECT 2553.160 82.870 2553.300 134.310 ;
        RECT 2553.160 82.730 2556.520 82.870 ;
        RECT 2556.380 2.400 2556.520 82.730 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 636.480 499.500 636.800 499.760 ;
        RECT 636.570 498.740 636.710 499.500 ;
        RECT 636.250 498.540 636.710 498.740 ;
        RECT 636.250 498.480 636.570 498.540 ;
        RECT 636.250 489.840 636.570 489.900 ;
        RECT 637.630 489.840 637.950 489.900 ;
        RECT 636.250 489.700 637.950 489.840 ;
        RECT 636.250 489.640 636.570 489.700 ;
        RECT 637.630 489.640 637.950 489.700 ;
        RECT 637.630 142.020 637.950 142.080 ;
        RECT 2574.230 142.020 2574.550 142.080 ;
        RECT 637.630 141.880 2574.550 142.020 ;
        RECT 637.630 141.820 637.950 141.880 ;
        RECT 2574.230 141.820 2574.550 141.880 ;
      LAYER via ;
        RECT 636.510 499.500 636.770 499.760 ;
        RECT 636.280 498.480 636.540 498.740 ;
        RECT 636.280 489.640 636.540 489.900 ;
        RECT 637.660 489.640 637.920 489.900 ;
        RECT 637.660 141.820 637.920 142.080 ;
        RECT 2574.260 141.820 2574.520 142.080 ;
      LAYER met2 ;
        RECT 636.530 500.000 636.810 504.000 ;
        RECT 636.570 499.790 636.710 500.000 ;
        RECT 636.510 499.470 636.770 499.790 ;
        RECT 636.280 498.450 636.540 498.770 ;
        RECT 636.340 489.930 636.480 498.450 ;
        RECT 636.280 489.610 636.540 489.930 ;
        RECT 637.660 489.610 637.920 489.930 ;
        RECT 637.720 142.110 637.860 489.610 ;
        RECT 637.660 141.790 637.920 142.110 ;
        RECT 2574.260 141.790 2574.520 142.110 ;
        RECT 2574.320 16.730 2574.460 141.790 ;
        RECT 2573.860 16.590 2574.460 16.730 ;
        RECT 2573.860 2.400 2574.000 16.590 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 500.090 171.940 500.410 172.000 ;
        RECT 814.270 171.940 814.590 172.000 ;
        RECT 500.090 171.800 814.590 171.940 ;
        RECT 500.090 171.740 500.410 171.800 ;
        RECT 814.270 171.740 814.590 171.800 ;
      LAYER via ;
        RECT 500.120 171.740 500.380 172.000 ;
        RECT 814.300 171.740 814.560 172.000 ;
      LAYER met2 ;
        RECT 499.910 500.000 500.190 504.000 ;
        RECT 499.950 499.815 500.090 500.000 ;
        RECT 499.880 499.445 500.160 499.815 ;
        RECT 500.110 498.595 500.390 498.965 ;
        RECT 500.180 172.030 500.320 498.595 ;
        RECT 500.120 171.710 500.380 172.030 ;
        RECT 814.300 171.710 814.560 172.030 ;
        RECT 814.360 82.870 814.500 171.710 ;
        RECT 814.360 82.730 818.640 82.870 ;
        RECT 818.500 2.400 818.640 82.730 ;
        RECT 818.290 -4.800 818.850 2.400 ;
      LAYER via2 ;
        RECT 499.880 499.490 500.160 499.770 ;
        RECT 500.110 498.640 500.390 498.920 ;
      LAYER met3 ;
        RECT 499.855 499.465 500.185 499.795 ;
        RECT 499.870 498.945 500.170 499.465 ;
        RECT 499.870 498.630 500.415 498.945 ;
        RECT 500.085 498.615 500.415 498.630 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 637.860 499.500 638.180 499.760 ;
        RECT 637.950 498.060 638.090 499.500 ;
        RECT 637.950 497.860 638.410 498.060 ;
        RECT 638.090 497.800 638.410 497.860 ;
        RECT 638.090 141.680 638.410 141.740 ;
        RECT 2587.570 141.680 2587.890 141.740 ;
        RECT 638.090 141.540 2587.890 141.680 ;
        RECT 638.090 141.480 638.410 141.540 ;
        RECT 2587.570 141.480 2587.890 141.540 ;
      LAYER via ;
        RECT 637.890 499.500 638.150 499.760 ;
        RECT 638.120 497.800 638.380 498.060 ;
        RECT 638.120 141.480 638.380 141.740 ;
        RECT 2587.600 141.480 2587.860 141.740 ;
      LAYER met2 ;
        RECT 637.910 500.000 638.190 504.000 ;
        RECT 637.950 499.790 638.090 500.000 ;
        RECT 637.890 499.470 638.150 499.790 ;
        RECT 638.120 497.770 638.380 498.090 ;
        RECT 638.180 141.770 638.320 497.770 ;
        RECT 638.120 141.450 638.380 141.770 ;
        RECT 2587.600 141.450 2587.860 141.770 ;
        RECT 2587.660 82.870 2587.800 141.450 ;
        RECT 2587.660 82.730 2589.640 82.870 ;
        RECT 2589.500 1.770 2589.640 82.730 ;
        RECT 2591.590 1.770 2592.150 2.400 ;
        RECT 2589.500 1.630 2592.150 1.770 ;
        RECT 2591.590 -4.800 2592.150 1.630 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 639.240 498.820 639.560 499.080 ;
        RECT 638.550 497.320 638.870 497.380 ;
        RECT 639.330 497.320 639.470 498.820 ;
        RECT 638.550 497.180 639.470 497.320 ;
        RECT 638.550 497.120 638.870 497.180 ;
        RECT 638.550 410.620 638.870 410.680 ;
        RECT 2608.270 410.620 2608.590 410.680 ;
        RECT 638.550 410.480 2608.590 410.620 ;
        RECT 638.550 410.420 638.870 410.480 ;
        RECT 2608.270 410.420 2608.590 410.480 ;
      LAYER via ;
        RECT 639.270 498.820 639.530 499.080 ;
        RECT 638.580 497.120 638.840 497.380 ;
        RECT 638.580 410.420 638.840 410.680 ;
        RECT 2608.300 410.420 2608.560 410.680 ;
      LAYER met2 ;
        RECT 639.290 500.000 639.570 504.000 ;
        RECT 639.330 499.110 639.470 500.000 ;
        RECT 639.270 498.790 639.530 499.110 ;
        RECT 638.580 497.090 638.840 497.410 ;
        RECT 638.640 410.710 638.780 497.090 ;
        RECT 638.580 410.390 638.840 410.710 ;
        RECT 2608.300 410.390 2608.560 410.710 ;
        RECT 2608.360 1.770 2608.500 410.390 ;
        RECT 2609.070 1.770 2609.630 2.400 ;
        RECT 2608.360 1.630 2609.630 1.770 ;
        RECT 2609.070 -4.800 2609.630 1.630 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.670 500.000 640.950 504.000 ;
        RECT 640.710 498.850 640.850 500.000 ;
        RECT 640.480 498.710 640.850 498.850 ;
        RECT 640.480 494.885 640.620 498.710 ;
        RECT 640.410 494.515 640.690 494.885 ;
        RECT 2622.090 141.595 2622.370 141.965 ;
        RECT 2622.160 82.870 2622.300 141.595 ;
        RECT 2622.160 82.730 2627.360 82.870 ;
        RECT 2627.220 2.400 2627.360 82.730 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
      LAYER via2 ;
        RECT 640.410 494.560 640.690 494.840 ;
        RECT 2622.090 141.640 2622.370 141.920 ;
      LAYER met3 ;
        RECT 635.990 494.850 636.370 494.860 ;
        RECT 640.385 494.850 640.715 494.865 ;
        RECT 635.990 494.550 640.715 494.850 ;
        RECT 635.990 494.540 636.370 494.550 ;
        RECT 640.385 494.535 640.715 494.550 ;
        RECT 635.990 141.930 636.370 141.940 ;
        RECT 2622.065 141.930 2622.395 141.945 ;
        RECT 635.990 141.630 2622.395 141.930 ;
        RECT 635.990 141.620 636.370 141.630 ;
        RECT 2622.065 141.615 2622.395 141.630 ;
      LAYER via3 ;
        RECT 636.020 494.540 636.340 494.860 ;
        RECT 636.020 141.620 636.340 141.940 ;
      LAYER met4 ;
        RECT 636.015 494.535 636.345 494.865 ;
        RECT 636.030 141.945 636.330 494.535 ;
        RECT 636.015 141.615 636.345 141.945 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 642.090 499.900 645.910 500.040 ;
        RECT 642.090 499.760 642.230 499.900 ;
        RECT 642.000 499.500 642.320 499.760 ;
        RECT 645.770 497.660 645.910 499.900 ;
        RECT 646.370 497.660 646.690 497.720 ;
        RECT 645.770 497.520 646.690 497.660 ;
        RECT 646.370 497.460 646.690 497.520 ;
        RECT 644.990 453.800 645.310 453.860 ;
        RECT 647.750 453.800 648.070 453.860 ;
        RECT 644.990 453.660 648.070 453.800 ;
        RECT 644.990 453.600 645.310 453.660 ;
        RECT 647.750 453.600 648.070 453.660 ;
        RECT 644.990 141.340 645.310 141.400 ;
        RECT 2642.770 141.340 2643.090 141.400 ;
        RECT 644.990 141.200 2643.090 141.340 ;
        RECT 644.990 141.140 645.310 141.200 ;
        RECT 2642.770 141.140 2643.090 141.200 ;
      LAYER via ;
        RECT 642.030 499.500 642.290 499.760 ;
        RECT 646.400 497.460 646.660 497.720 ;
        RECT 645.020 453.600 645.280 453.860 ;
        RECT 647.780 453.600 648.040 453.860 ;
        RECT 645.020 141.140 645.280 141.400 ;
        RECT 2642.800 141.140 2643.060 141.400 ;
      LAYER met2 ;
        RECT 642.050 500.000 642.330 504.000 ;
        RECT 642.090 499.790 642.230 500.000 ;
        RECT 642.030 499.470 642.290 499.790 ;
        RECT 646.400 497.430 646.660 497.750 ;
        RECT 646.460 476.170 646.600 497.430 ;
        RECT 646.460 476.030 647.980 476.170 ;
        RECT 647.840 453.890 647.980 476.030 ;
        RECT 645.020 453.570 645.280 453.890 ;
        RECT 647.780 453.570 648.040 453.890 ;
        RECT 645.080 141.430 645.220 453.570 ;
        RECT 645.020 141.110 645.280 141.430 ;
        RECT 2642.800 141.110 2643.060 141.430 ;
        RECT 2642.860 1.770 2643.000 141.110 ;
        RECT 2644.950 1.770 2645.510 2.400 ;
        RECT 2642.860 1.630 2645.510 1.770 ;
        RECT 2644.950 -4.800 2645.510 1.630 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 643.380 499.500 643.700 499.760 ;
        RECT 643.470 497.320 643.610 499.500 ;
        RECT 644.990 497.320 645.310 497.380 ;
        RECT 643.470 497.180 645.310 497.320 ;
        RECT 644.990 497.120 645.310 497.180 ;
        RECT 644.990 473.520 645.310 473.580 ;
        RECT 646.370 473.520 646.690 473.580 ;
        RECT 644.990 473.380 646.690 473.520 ;
        RECT 644.990 473.320 645.310 473.380 ;
        RECT 646.370 473.320 646.690 473.380 ;
        RECT 645.910 149.160 646.230 149.220 ;
        RECT 2656.570 149.160 2656.890 149.220 ;
        RECT 645.910 149.020 2656.890 149.160 ;
        RECT 645.910 148.960 646.230 149.020 ;
        RECT 2656.570 148.960 2656.890 149.020 ;
        RECT 2656.570 17.580 2656.890 17.640 ;
        RECT 2660.710 17.580 2661.030 17.640 ;
        RECT 2656.570 17.440 2661.030 17.580 ;
        RECT 2656.570 17.380 2656.890 17.440 ;
        RECT 2660.710 17.380 2661.030 17.440 ;
      LAYER via ;
        RECT 643.410 499.500 643.670 499.760 ;
        RECT 645.020 497.120 645.280 497.380 ;
        RECT 645.020 473.320 645.280 473.580 ;
        RECT 646.400 473.320 646.660 473.580 ;
        RECT 645.940 148.960 646.200 149.220 ;
        RECT 2656.600 148.960 2656.860 149.220 ;
        RECT 2656.600 17.380 2656.860 17.640 ;
        RECT 2660.740 17.380 2661.000 17.640 ;
      LAYER met2 ;
        RECT 643.430 500.000 643.710 504.000 ;
        RECT 643.470 499.790 643.610 500.000 ;
        RECT 643.410 499.470 643.670 499.790 ;
        RECT 645.020 497.090 645.280 497.410 ;
        RECT 645.080 473.610 645.220 497.090 ;
        RECT 645.020 473.290 645.280 473.610 ;
        RECT 646.400 473.290 646.660 473.610 ;
        RECT 646.460 448.570 646.600 473.290 ;
        RECT 646.000 448.430 646.600 448.570 ;
        RECT 646.000 149.250 646.140 448.430 ;
        RECT 645.940 148.930 646.200 149.250 ;
        RECT 2656.600 148.930 2656.860 149.250 ;
        RECT 2656.660 17.670 2656.800 148.930 ;
        RECT 2656.600 17.350 2656.860 17.670 ;
        RECT 2660.740 17.350 2661.000 17.670 ;
        RECT 2660.800 1.770 2660.940 17.350 ;
        RECT 2662.430 1.770 2662.990 2.400 ;
        RECT 2660.800 1.630 2662.990 1.770 ;
        RECT 2662.430 -4.800 2662.990 1.630 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 644.760 499.700 645.080 499.760 ;
        RECT 644.620 499.500 645.080 499.700 ;
        RECT 644.620 499.080 644.760 499.500 ;
        RECT 644.530 498.820 644.850 499.080 ;
        RECT 645.450 148.820 645.770 148.880 ;
        RECT 2677.270 148.820 2677.590 148.880 ;
        RECT 645.450 148.680 2677.590 148.820 ;
        RECT 645.450 148.620 645.770 148.680 ;
        RECT 2677.270 148.620 2677.590 148.680 ;
      LAYER via ;
        RECT 644.790 499.500 645.050 499.760 ;
        RECT 644.560 498.820 644.820 499.080 ;
        RECT 645.480 148.620 645.740 148.880 ;
        RECT 2677.300 148.620 2677.560 148.880 ;
      LAYER met2 ;
        RECT 644.810 500.000 645.090 504.000 ;
        RECT 644.850 499.790 644.990 500.000 ;
        RECT 644.790 499.470 645.050 499.790 ;
        RECT 644.560 498.790 644.820 499.110 ;
        RECT 644.620 473.010 644.760 498.790 ;
        RECT 644.620 472.870 645.680 473.010 ;
        RECT 645.540 148.910 645.680 472.870 ;
        RECT 645.480 148.590 645.740 148.910 ;
        RECT 2677.300 148.590 2677.560 148.910 ;
        RECT 2677.360 82.870 2677.500 148.590 ;
        RECT 2677.360 82.730 2680.720 82.870 ;
        RECT 2680.580 2.400 2680.720 82.730 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.190 500.000 646.470 504.000 ;
        RECT 646.230 499.815 646.370 500.000 ;
        RECT 646.160 499.445 646.440 499.815 ;
        RECT 2697.990 140.915 2698.270 141.285 ;
        RECT 2698.060 2.400 2698.200 140.915 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
      LAYER via2 ;
        RECT 646.160 499.490 646.440 499.770 ;
        RECT 2697.990 140.960 2698.270 141.240 ;
      LAYER met3 ;
        RECT 646.135 499.620 646.465 499.795 ;
        RECT 646.110 499.610 646.490 499.620 ;
        RECT 646.110 499.310 646.750 499.610 ;
        RECT 646.110 499.300 646.490 499.310 ;
        RECT 646.110 141.250 646.490 141.260 ;
        RECT 2697.965 141.250 2698.295 141.265 ;
        RECT 646.110 140.950 2698.295 141.250 ;
        RECT 646.110 140.940 646.490 140.950 ;
        RECT 2697.965 140.935 2698.295 140.950 ;
      LAYER via3 ;
        RECT 646.140 499.300 646.460 499.620 ;
        RECT 646.140 140.940 646.460 141.260 ;
      LAYER met4 ;
        RECT 646.135 499.295 646.465 499.625 ;
        RECT 646.150 141.265 646.450 499.295 ;
        RECT 646.135 140.935 646.465 141.265 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 647.520 499.360 647.840 499.420 ;
        RECT 647.520 499.160 647.980 499.360 ;
        RECT 647.840 498.060 647.980 499.160 ;
        RECT 647.750 497.800 648.070 498.060 ;
      LAYER via ;
        RECT 647.550 499.160 647.810 499.420 ;
        RECT 647.780 497.800 648.040 498.060 ;
      LAYER met2 ;
        RECT 647.570 500.000 647.850 504.000 ;
        RECT 647.610 499.450 647.750 500.000 ;
        RECT 647.550 499.130 647.810 499.450 ;
        RECT 647.780 497.770 648.040 498.090 ;
        RECT 647.840 487.405 647.980 497.770 ;
        RECT 647.770 487.035 648.050 487.405 ;
        RECT 2711.790 176.955 2712.070 177.325 ;
        RECT 2711.860 82.870 2712.000 176.955 ;
        RECT 2711.860 82.730 2713.840 82.870 ;
        RECT 2713.700 1.770 2713.840 82.730 ;
        RECT 2715.790 1.770 2716.350 2.400 ;
        RECT 2713.700 1.630 2716.350 1.770 ;
        RECT 2715.790 -4.800 2716.350 1.630 ;
      LAYER via2 ;
        RECT 647.770 487.080 648.050 487.360 ;
        RECT 2711.790 177.000 2712.070 177.280 ;
      LAYER met3 ;
        RECT 645.190 487.370 645.570 487.380 ;
        RECT 647.745 487.370 648.075 487.385 ;
        RECT 645.190 487.070 648.075 487.370 ;
        RECT 645.190 487.060 645.570 487.070 ;
        RECT 647.745 487.055 648.075 487.070 ;
        RECT 645.190 177.290 645.570 177.300 ;
        RECT 2711.765 177.290 2712.095 177.305 ;
        RECT 645.190 176.990 2712.095 177.290 ;
        RECT 645.190 176.980 645.570 176.990 ;
        RECT 2711.765 176.975 2712.095 176.990 ;
      LAYER via3 ;
        RECT 645.220 487.060 645.540 487.380 ;
        RECT 645.220 176.980 645.540 177.300 ;
      LAYER met4 ;
        RECT 645.215 487.055 645.545 487.385 ;
        RECT 645.230 177.305 645.530 487.055 ;
        RECT 645.215 176.975 645.545 177.305 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 648.900 499.160 649.220 499.420 ;
        RECT 648.990 498.000 649.130 499.160 ;
        RECT 649.590 498.000 649.910 498.060 ;
        RECT 648.990 497.860 649.910 498.000 ;
        RECT 649.590 497.800 649.910 497.860 ;
        RECT 651.890 148.480 652.210 148.540 ;
        RECT 2732.470 148.480 2732.790 148.540 ;
        RECT 651.890 148.340 2732.790 148.480 ;
        RECT 651.890 148.280 652.210 148.340 ;
        RECT 2732.470 148.280 2732.790 148.340 ;
      LAYER via ;
        RECT 648.930 499.160 649.190 499.420 ;
        RECT 649.620 497.800 649.880 498.060 ;
        RECT 651.920 148.280 652.180 148.540 ;
        RECT 2732.500 148.280 2732.760 148.540 ;
      LAYER met2 ;
        RECT 648.950 500.000 649.230 504.000 ;
        RECT 648.990 499.450 649.130 500.000 ;
        RECT 648.930 499.130 649.190 499.450 ;
        RECT 649.620 497.770 649.880 498.090 ;
        RECT 649.680 475.165 649.820 497.770 ;
        RECT 649.610 474.795 649.890 475.165 ;
        RECT 651.910 472.075 652.190 472.445 ;
        RECT 651.980 148.570 652.120 472.075 ;
        RECT 651.920 148.250 652.180 148.570 ;
        RECT 2732.500 148.250 2732.760 148.570 ;
        RECT 2732.560 1.770 2732.700 148.250 ;
        RECT 2733.270 1.770 2733.830 2.400 ;
        RECT 2732.560 1.630 2733.830 1.770 ;
        RECT 2733.270 -4.800 2733.830 1.630 ;
      LAYER via2 ;
        RECT 649.610 474.840 649.890 475.120 ;
        RECT 651.910 472.120 652.190 472.400 ;
      LAYER met3 ;
        RECT 649.585 475.130 649.915 475.145 ;
        RECT 649.585 474.830 651.050 475.130 ;
        RECT 649.585 474.815 649.915 474.830 ;
        RECT 650.750 472.410 651.050 474.830 ;
        RECT 651.885 472.410 652.215 472.425 ;
        RECT 650.750 472.110 652.215 472.410 ;
        RECT 651.885 472.095 652.215 472.110 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 651.430 148.140 651.750 148.200 ;
        RECT 2746.270 148.140 2746.590 148.200 ;
        RECT 651.430 148.000 2746.590 148.140 ;
        RECT 651.430 147.940 651.750 148.000 ;
        RECT 2746.270 147.940 2746.590 148.000 ;
      LAYER via ;
        RECT 651.460 147.940 651.720 148.200 ;
        RECT 2746.300 147.940 2746.560 148.200 ;
      LAYER met2 ;
        RECT 650.330 500.000 650.610 504.000 ;
        RECT 650.370 499.815 650.510 500.000 ;
        RECT 650.300 499.445 650.580 499.815 ;
        RECT 651.450 497.915 651.730 498.285 ;
        RECT 651.520 148.230 651.660 497.915 ;
        RECT 651.460 147.910 651.720 148.230 ;
        RECT 2746.300 147.910 2746.560 148.230 ;
        RECT 2746.360 82.870 2746.500 147.910 ;
        RECT 2746.360 82.730 2751.560 82.870 ;
        RECT 2751.420 2.400 2751.560 82.730 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
      LAYER via2 ;
        RECT 650.300 499.490 650.580 499.770 ;
        RECT 651.450 497.960 651.730 498.240 ;
      LAYER met3 ;
        RECT 650.275 499.780 650.605 499.795 ;
        RECT 650.275 499.610 650.820 499.780 ;
        RECT 650.275 499.465 651.970 499.610 ;
        RECT 650.520 499.310 651.970 499.465 ;
        RECT 651.670 498.265 651.970 499.310 ;
        RECT 651.425 497.950 651.970 498.265 ;
        RECT 651.425 497.935 651.755 497.950 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 500.550 177.720 500.870 177.780 ;
        RECT 834.970 177.720 835.290 177.780 ;
        RECT 500.550 177.580 835.290 177.720 ;
        RECT 500.550 177.520 500.870 177.580 ;
        RECT 834.970 177.520 835.290 177.580 ;
      LAYER via ;
        RECT 500.580 177.520 500.840 177.780 ;
        RECT 835.000 177.520 835.260 177.780 ;
      LAYER met2 ;
        RECT 501.290 500.000 501.570 504.000 ;
        RECT 501.330 498.680 501.470 500.000 ;
        RECT 501.100 498.540 501.470 498.680 ;
        RECT 501.100 498.340 501.240 498.540 ;
        RECT 500.640 498.200 501.240 498.340 ;
        RECT 500.640 177.810 500.780 498.200 ;
        RECT 500.580 177.490 500.840 177.810 ;
        RECT 835.000 177.490 835.260 177.810 ;
        RECT 835.060 82.870 835.200 177.490 ;
        RECT 835.060 82.730 836.120 82.870 ;
        RECT 835.980 2.400 836.120 82.730 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 651.890 472.840 652.210 472.900 ;
        RECT 652.810 472.840 653.130 472.900 ;
        RECT 651.890 472.700 653.130 472.840 ;
        RECT 651.890 472.640 652.210 472.700 ;
        RECT 652.810 472.640 653.130 472.700 ;
        RECT 652.810 176.020 653.130 176.080 ;
        RECT 2766.970 176.020 2767.290 176.080 ;
        RECT 652.810 175.880 2767.290 176.020 ;
        RECT 652.810 175.820 653.130 175.880 ;
        RECT 2766.970 175.820 2767.290 175.880 ;
      LAYER via ;
        RECT 651.920 472.640 652.180 472.900 ;
        RECT 652.840 472.640 653.100 472.900 ;
        RECT 652.840 175.820 653.100 176.080 ;
        RECT 2767.000 175.820 2767.260 176.080 ;
      LAYER met2 ;
        RECT 651.710 500.000 651.990 504.000 ;
        RECT 651.750 498.850 651.890 500.000 ;
        RECT 651.750 498.710 652.120 498.850 ;
        RECT 651.980 472.930 652.120 498.710 ;
        RECT 651.920 472.610 652.180 472.930 ;
        RECT 652.840 472.610 653.100 472.930 ;
        RECT 652.900 176.110 653.040 472.610 ;
        RECT 652.840 175.790 653.100 176.110 ;
        RECT 2767.000 175.790 2767.260 176.110 ;
        RECT 2767.060 82.870 2767.200 175.790 ;
        RECT 2767.060 82.730 2769.040 82.870 ;
        RECT 2768.900 2.400 2769.040 82.730 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 653.040 499.500 653.360 499.760 ;
        RECT 653.130 498.000 653.270 499.500 ;
        RECT 653.130 497.860 654.190 498.000 ;
        RECT 654.050 497.720 654.190 497.860 ;
        RECT 654.050 497.520 654.510 497.720 ;
        RECT 654.190 497.460 654.510 497.520 ;
        RECT 652.350 488.480 652.670 488.540 ;
        RECT 654.190 488.480 654.510 488.540 ;
        RECT 652.350 488.340 654.510 488.480 ;
        RECT 652.350 488.280 652.670 488.340 ;
        RECT 654.190 488.280 654.510 488.340 ;
        RECT 652.350 155.280 652.670 155.340 ;
        RECT 2780.770 155.280 2781.090 155.340 ;
        RECT 652.350 155.140 2781.090 155.280 ;
        RECT 652.350 155.080 652.670 155.140 ;
        RECT 2780.770 155.080 2781.090 155.140 ;
        RECT 2780.770 17.580 2781.090 17.640 ;
        RECT 2784.910 17.580 2785.230 17.640 ;
        RECT 2780.770 17.440 2785.230 17.580 ;
        RECT 2780.770 17.380 2781.090 17.440 ;
        RECT 2784.910 17.380 2785.230 17.440 ;
      LAYER via ;
        RECT 653.070 499.500 653.330 499.760 ;
        RECT 654.220 497.460 654.480 497.720 ;
        RECT 652.380 488.280 652.640 488.540 ;
        RECT 654.220 488.280 654.480 488.540 ;
        RECT 652.380 155.080 652.640 155.340 ;
        RECT 2780.800 155.080 2781.060 155.340 ;
        RECT 2780.800 17.380 2781.060 17.640 ;
        RECT 2784.940 17.380 2785.200 17.640 ;
      LAYER met2 ;
        RECT 653.090 500.000 653.370 504.000 ;
        RECT 653.130 499.790 653.270 500.000 ;
        RECT 653.070 499.470 653.330 499.790 ;
        RECT 654.220 497.430 654.480 497.750 ;
        RECT 654.280 488.570 654.420 497.430 ;
        RECT 652.380 488.250 652.640 488.570 ;
        RECT 654.220 488.250 654.480 488.570 ;
        RECT 652.440 155.370 652.580 488.250 ;
        RECT 652.380 155.050 652.640 155.370 ;
        RECT 2780.800 155.050 2781.060 155.370 ;
        RECT 2780.860 17.670 2781.000 155.050 ;
        RECT 2780.800 17.350 2781.060 17.670 ;
        RECT 2784.940 17.350 2785.200 17.670 ;
        RECT 2785.000 1.770 2785.140 17.350 ;
        RECT 2786.630 1.770 2787.190 2.400 ;
        RECT 2785.000 1.630 2787.190 1.770 ;
        RECT 2786.630 -4.800 2787.190 1.630 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.470 500.000 654.750 504.000 ;
        RECT 654.510 498.680 654.650 500.000 ;
        RECT 654.510 498.540 654.880 498.680 ;
        RECT 654.740 491.485 654.880 498.540 ;
        RECT 654.670 491.115 654.950 491.485 ;
        RECT 2801.490 176.275 2801.770 176.645 ;
        RECT 2801.560 82.870 2801.700 176.275 ;
        RECT 2801.560 82.730 2802.160 82.870 ;
        RECT 2802.020 1.770 2802.160 82.730 ;
        RECT 2804.110 1.770 2804.670 2.400 ;
        RECT 2802.020 1.630 2804.670 1.770 ;
        RECT 2804.110 -4.800 2804.670 1.630 ;
      LAYER via2 ;
        RECT 654.670 491.160 654.950 491.440 ;
        RECT 2801.490 176.320 2801.770 176.600 ;
      LAYER met3 ;
        RECT 651.630 491.450 652.010 491.460 ;
        RECT 654.645 491.450 654.975 491.465 ;
        RECT 651.630 491.150 654.975 491.450 ;
        RECT 651.630 491.140 652.010 491.150 ;
        RECT 654.645 491.135 654.975 491.150 ;
        RECT 651.630 176.610 652.010 176.620 ;
        RECT 2801.465 176.610 2801.795 176.625 ;
        RECT 651.630 176.310 2801.795 176.610 ;
        RECT 651.630 176.300 652.010 176.310 ;
        RECT 2801.465 176.295 2801.795 176.310 ;
      LAYER via3 ;
        RECT 651.660 491.140 651.980 491.460 ;
        RECT 651.660 176.300 651.980 176.620 ;
      LAYER met4 ;
        RECT 651.655 491.135 651.985 491.465 ;
        RECT 651.670 176.625 651.970 491.135 ;
        RECT 651.655 176.295 651.985 176.625 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.030 472.500 656.350 472.560 ;
        RECT 658.790 472.500 659.110 472.560 ;
        RECT 656.030 472.360 659.110 472.500 ;
        RECT 656.030 472.300 656.350 472.360 ;
        RECT 658.790 472.300 659.110 472.360 ;
        RECT 658.790 100.200 659.110 100.260 ;
        RECT 2822.170 100.200 2822.490 100.260 ;
        RECT 658.790 100.060 2822.490 100.200 ;
        RECT 658.790 100.000 659.110 100.060 ;
        RECT 2822.170 100.000 2822.490 100.060 ;
      LAYER via ;
        RECT 656.060 472.300 656.320 472.560 ;
        RECT 658.820 472.300 659.080 472.560 ;
        RECT 658.820 100.000 659.080 100.260 ;
        RECT 2822.200 100.000 2822.460 100.260 ;
      LAYER met2 ;
        RECT 655.850 500.000 656.130 504.000 ;
        RECT 655.890 498.680 656.030 500.000 ;
        RECT 655.890 498.540 656.260 498.680 ;
        RECT 656.120 472.590 656.260 498.540 ;
        RECT 656.060 472.270 656.320 472.590 ;
        RECT 658.820 472.270 659.080 472.590 ;
        RECT 658.880 100.290 659.020 472.270 ;
        RECT 658.820 99.970 659.080 100.290 ;
        RECT 2822.200 99.970 2822.460 100.290 ;
        RECT 2822.260 2.400 2822.400 99.970 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.950 489.840 657.270 489.900 ;
        RECT 658.790 489.840 659.110 489.900 ;
        RECT 656.950 489.700 659.110 489.840 ;
        RECT 656.950 489.640 657.270 489.700 ;
        RECT 658.790 489.640 659.110 489.700 ;
        RECT 659.250 162.080 659.570 162.140 ;
        RECT 2835.970 162.080 2836.290 162.140 ;
        RECT 659.250 161.940 2836.290 162.080 ;
        RECT 659.250 161.880 659.570 161.940 ;
        RECT 2835.970 161.880 2836.290 161.940 ;
      LAYER via ;
        RECT 656.980 489.640 657.240 489.900 ;
        RECT 658.820 489.640 659.080 489.900 ;
        RECT 659.280 161.880 659.540 162.140 ;
        RECT 2836.000 161.880 2836.260 162.140 ;
      LAYER met2 ;
        RECT 657.230 500.000 657.510 504.000 ;
        RECT 657.270 498.680 657.410 500.000 ;
        RECT 657.040 498.540 657.410 498.680 ;
        RECT 657.040 489.930 657.180 498.540 ;
        RECT 656.980 489.610 657.240 489.930 ;
        RECT 658.820 489.610 659.080 489.930 ;
        RECT 658.880 473.010 659.020 489.610 ;
        RECT 658.880 472.870 659.480 473.010 ;
        RECT 659.340 162.170 659.480 472.870 ;
        RECT 659.280 161.850 659.540 162.170 ;
        RECT 2836.000 161.850 2836.260 162.170 ;
        RECT 2836.060 82.870 2836.200 161.850 ;
        RECT 2836.060 82.730 2838.040 82.870 ;
        RECT 2837.900 1.770 2838.040 82.730 ;
        RECT 2839.990 1.770 2840.550 2.400 ;
        RECT 2837.900 1.630 2840.550 1.770 ;
        RECT 2839.990 -4.800 2840.550 1.630 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 658.560 499.360 658.880 499.420 ;
        RECT 658.420 499.160 658.880 499.360 ;
        RECT 658.420 497.380 658.560 499.160 ;
        RECT 658.330 497.120 658.650 497.380 ;
        RECT 658.330 99.860 658.650 99.920 ;
        RECT 2856.670 99.860 2856.990 99.920 ;
        RECT 658.330 99.720 2856.990 99.860 ;
        RECT 658.330 99.660 658.650 99.720 ;
        RECT 2856.670 99.660 2856.990 99.720 ;
      LAYER via ;
        RECT 658.590 499.160 658.850 499.420 ;
        RECT 658.360 497.120 658.620 497.380 ;
        RECT 658.360 99.660 658.620 99.920 ;
        RECT 2856.700 99.660 2856.960 99.920 ;
      LAYER met2 ;
        RECT 658.610 500.000 658.890 504.000 ;
        RECT 658.650 499.450 658.790 500.000 ;
        RECT 658.590 499.130 658.850 499.450 ;
        RECT 658.360 497.090 658.620 497.410 ;
        RECT 658.420 99.950 658.560 497.090 ;
        RECT 658.360 99.630 658.620 99.950 ;
        RECT 2856.700 99.630 2856.960 99.950 ;
        RECT 2856.760 1.770 2856.900 99.630 ;
        RECT 2857.470 1.770 2858.030 2.400 ;
        RECT 2856.760 1.630 2858.030 1.770 ;
        RECT 2857.470 -4.800 2858.030 1.630 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.990 500.000 660.270 504.000 ;
        RECT 660.030 499.645 660.170 500.000 ;
        RECT 659.960 499.275 660.240 499.645 ;
        RECT 2870.490 175.595 2870.770 175.965 ;
        RECT 2870.560 82.870 2870.700 175.595 ;
        RECT 2870.560 82.730 2875.760 82.870 ;
        RECT 2875.620 2.400 2875.760 82.730 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
      LAYER via2 ;
        RECT 659.960 499.320 660.240 499.600 ;
        RECT 2870.490 175.640 2870.770 175.920 ;
      LAYER met3 ;
        RECT 659.935 499.620 660.265 499.625 ;
        RECT 659.910 499.610 660.290 499.620 ;
        RECT 659.910 499.310 660.720 499.610 ;
        RECT 659.910 499.300 660.290 499.310 ;
        RECT 659.935 499.295 660.265 499.300 ;
        RECT 657.150 175.930 657.530 175.940 ;
        RECT 2870.465 175.930 2870.795 175.945 ;
        RECT 657.150 175.630 2870.795 175.930 ;
        RECT 657.150 175.620 657.530 175.630 ;
        RECT 2870.465 175.615 2870.795 175.630 ;
      LAYER via3 ;
        RECT 659.940 499.300 660.260 499.620 ;
        RECT 657.180 175.620 657.500 175.940 ;
      LAYER met4 ;
        RECT 659.935 499.610 660.265 499.625 ;
        RECT 657.190 499.310 660.265 499.610 ;
        RECT 657.190 175.945 657.490 499.310 ;
        RECT 659.935 499.295 660.265 499.310 ;
        RECT 657.175 175.615 657.505 175.945 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.370 500.000 661.650 504.000 ;
        RECT 661.410 499.645 661.550 500.000 ;
        RECT 661.340 499.275 661.620 499.645 ;
        RECT 2891.190 99.435 2891.470 99.805 ;
        RECT 2891.260 82.870 2891.400 99.435 ;
        RECT 2891.260 82.730 2893.240 82.870 ;
        RECT 2893.100 2.400 2893.240 82.730 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
      LAYER via2 ;
        RECT 661.340 499.320 661.620 499.600 ;
        RECT 2891.190 99.480 2891.470 99.760 ;
      LAYER met3 ;
        RECT 661.315 499.295 661.645 499.625 ;
        RECT 659.910 498.930 660.290 498.940 ;
        RECT 661.330 498.930 661.630 499.295 ;
        RECT 659.910 498.630 661.630 498.930 ;
        RECT 659.910 498.620 660.290 498.630 ;
        RECT 658.990 99.770 659.370 99.780 ;
        RECT 2891.165 99.770 2891.495 99.785 ;
        RECT 658.990 99.470 2891.495 99.770 ;
        RECT 658.990 99.460 659.370 99.470 ;
        RECT 2891.165 99.455 2891.495 99.470 ;
      LAYER via3 ;
        RECT 659.940 498.620 660.260 498.940 ;
        RECT 659.020 99.460 659.340 99.780 ;
      LAYER met4 ;
        RECT 659.935 498.930 660.265 498.945 ;
        RECT 659.030 498.630 660.265 498.930 ;
        RECT 659.030 99.785 659.330 498.630 ;
        RECT 659.935 498.615 660.265 498.630 ;
        RECT 659.015 99.455 659.345 99.785 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.670 500.000 502.950 504.000 ;
        RECT 502.710 498.340 502.850 500.000 ;
        RECT 502.480 498.200 502.850 498.340 ;
        RECT 502.480 492.165 502.620 498.200 ;
        RECT 502.410 491.795 502.690 492.165 ;
        RECT 848.790 178.315 849.070 178.685 ;
        RECT 848.860 82.870 849.000 178.315 ;
        RECT 848.860 82.730 851.760 82.870 ;
        RECT 851.620 1.770 851.760 82.730 ;
        RECT 853.710 1.770 854.270 2.400 ;
        RECT 851.620 1.630 854.270 1.770 ;
        RECT 853.710 -4.800 854.270 1.630 ;
      LAYER via2 ;
        RECT 502.410 491.840 502.690 492.120 ;
        RECT 848.790 178.360 849.070 178.640 ;
      LAYER met3 ;
        RECT 499.830 492.130 500.210 492.140 ;
        RECT 502.385 492.130 502.715 492.145 ;
        RECT 499.830 491.830 502.715 492.130 ;
        RECT 499.830 491.820 500.210 491.830 ;
        RECT 502.385 491.815 502.715 491.830 ;
        RECT 499.830 178.650 500.210 178.660 ;
        RECT 848.765 178.650 849.095 178.665 ;
        RECT 499.830 178.350 849.095 178.650 ;
        RECT 499.830 178.340 500.210 178.350 ;
        RECT 848.765 178.335 849.095 178.350 ;
      LAYER via3 ;
        RECT 499.860 491.820 500.180 492.140 ;
        RECT 499.860 178.340 500.180 178.660 ;
      LAYER met4 ;
        RECT 499.855 491.815 500.185 492.145 ;
        RECT 499.870 178.665 500.170 491.815 ;
        RECT 499.855 178.335 500.185 178.665 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.000 499.500 504.320 499.760 ;
        RECT 504.090 498.060 504.230 499.500 ;
        RECT 504.090 497.860 504.550 498.060 ;
        RECT 504.230 497.800 504.550 497.860 ;
        RECT 504.230 491.540 504.550 491.600 ;
        RECT 507.910 491.540 508.230 491.600 ;
        RECT 504.230 491.400 508.230 491.540 ;
        RECT 504.230 491.340 504.550 491.400 ;
        RECT 507.910 491.340 508.230 491.400 ;
        RECT 507.450 177.380 507.770 177.440 ;
        RECT 869.470 177.380 869.790 177.440 ;
        RECT 507.450 177.240 869.790 177.380 ;
        RECT 507.450 177.180 507.770 177.240 ;
        RECT 869.470 177.180 869.790 177.240 ;
      LAYER via ;
        RECT 504.030 499.500 504.290 499.760 ;
        RECT 504.260 497.800 504.520 498.060 ;
        RECT 504.260 491.340 504.520 491.600 ;
        RECT 507.940 491.340 508.200 491.600 ;
        RECT 507.480 177.180 507.740 177.440 ;
        RECT 869.500 177.180 869.760 177.440 ;
      LAYER met2 ;
        RECT 504.050 500.000 504.330 504.000 ;
        RECT 504.090 499.790 504.230 500.000 ;
        RECT 504.030 499.470 504.290 499.790 ;
        RECT 504.260 497.770 504.520 498.090 ;
        RECT 504.320 491.630 504.460 497.770 ;
        RECT 504.260 491.310 504.520 491.630 ;
        RECT 507.940 491.310 508.200 491.630 ;
        RECT 508.000 472.330 508.140 491.310 ;
        RECT 507.540 472.190 508.140 472.330 ;
        RECT 507.540 177.470 507.680 472.190 ;
        RECT 507.480 177.150 507.740 177.470 ;
        RECT 869.500 177.150 869.760 177.470 ;
        RECT 869.560 1.770 869.700 177.150 ;
        RECT 871.190 1.770 871.750 2.400 ;
        RECT 869.560 1.630 871.750 1.770 ;
        RECT 871.190 -4.800 871.750 1.630 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 506.530 177.040 506.850 177.100 ;
        RECT 883.270 177.040 883.590 177.100 ;
        RECT 506.530 176.900 883.590 177.040 ;
        RECT 506.530 176.840 506.850 176.900 ;
        RECT 883.270 176.840 883.590 176.900 ;
        RECT 883.270 58.380 883.590 58.440 ;
        RECT 889.250 58.380 889.570 58.440 ;
        RECT 883.270 58.240 889.570 58.380 ;
        RECT 883.270 58.180 883.590 58.240 ;
        RECT 889.250 58.180 889.570 58.240 ;
      LAYER via ;
        RECT 506.560 176.840 506.820 177.100 ;
        RECT 883.300 176.840 883.560 177.100 ;
        RECT 883.300 58.180 883.560 58.440 ;
        RECT 889.280 58.180 889.540 58.440 ;
      LAYER met2 ;
        RECT 505.430 500.000 505.710 504.000 ;
        RECT 505.470 499.645 505.610 500.000 ;
        RECT 505.400 499.275 505.680 499.645 ;
        RECT 506.090 497.235 506.370 497.605 ;
        RECT 506.160 472.500 506.300 497.235 ;
        RECT 506.160 472.360 506.760 472.500 ;
        RECT 506.620 177.130 506.760 472.360 ;
        RECT 506.560 176.810 506.820 177.130 ;
        RECT 883.300 176.810 883.560 177.130 ;
        RECT 883.360 58.470 883.500 176.810 ;
        RECT 883.300 58.150 883.560 58.470 ;
        RECT 889.280 58.150 889.540 58.470 ;
        RECT 889.340 2.400 889.480 58.150 ;
        RECT 889.130 -4.800 889.690 2.400 ;
      LAYER via2 ;
        RECT 505.400 499.320 505.680 499.600 ;
        RECT 506.090 497.280 506.370 497.560 ;
      LAYER met3 ;
        RECT 505.375 499.295 505.705 499.625 ;
        RECT 505.390 497.570 505.690 499.295 ;
        RECT 506.065 497.570 506.395 497.585 ;
        RECT 505.390 497.270 506.395 497.570 ;
        RECT 506.065 497.255 506.395 497.270 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 506.990 176.700 507.310 176.760 ;
        RECT 903.970 176.700 904.290 176.760 ;
        RECT 506.990 176.560 904.290 176.700 ;
        RECT 506.990 176.500 507.310 176.560 ;
        RECT 903.970 176.500 904.290 176.560 ;
      LAYER via ;
        RECT 507.020 176.500 507.280 176.760 ;
        RECT 904.000 176.500 904.260 176.760 ;
      LAYER met2 ;
        RECT 506.810 500.000 507.090 504.000 ;
        RECT 506.850 498.340 506.990 500.000 ;
        RECT 506.850 498.200 507.220 498.340 ;
        RECT 507.080 176.790 507.220 498.200 ;
        RECT 507.020 176.470 507.280 176.790 ;
        RECT 904.000 176.470 904.260 176.790 ;
        RECT 904.060 82.870 904.200 176.470 ;
        RECT 904.060 82.730 905.120 82.870 ;
        RECT 904.980 1.770 905.120 82.730 ;
        RECT 907.070 1.770 907.630 2.400 ;
        RECT 904.980 1.630 907.630 1.770 ;
        RECT 907.070 -4.800 907.630 1.630 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 508.140 499.160 508.460 499.420 ;
        RECT 508.230 498.400 508.370 499.160 ;
        RECT 508.230 498.200 508.690 498.400 ;
        RECT 508.370 498.140 508.690 498.200 ;
        RECT 508.370 492.360 508.690 492.620 ;
        RECT 508.460 491.880 508.600 492.360 ;
        RECT 530.910 491.880 531.230 491.940 ;
        RECT 508.460 491.740 531.230 491.880 ;
        RECT 530.910 491.680 531.230 491.740 ;
        RECT 530.910 487.800 531.230 487.860 ;
        RECT 570.470 487.800 570.790 487.860 ;
        RECT 530.910 487.660 570.790 487.800 ;
        RECT 530.910 487.600 531.230 487.660 ;
        RECT 570.470 487.600 570.790 487.660 ;
        RECT 570.470 182.140 570.790 182.200 ;
        RECT 924.670 182.140 924.990 182.200 ;
        RECT 570.470 182.000 924.990 182.140 ;
        RECT 570.470 181.940 570.790 182.000 ;
        RECT 924.670 181.940 924.990 182.000 ;
      LAYER via ;
        RECT 508.170 499.160 508.430 499.420 ;
        RECT 508.400 498.140 508.660 498.400 ;
        RECT 508.400 492.360 508.660 492.620 ;
        RECT 530.940 491.680 531.200 491.940 ;
        RECT 530.940 487.600 531.200 487.860 ;
        RECT 570.500 487.600 570.760 487.860 ;
        RECT 570.500 181.940 570.760 182.200 ;
        RECT 924.700 181.940 924.960 182.200 ;
      LAYER met2 ;
        RECT 508.190 500.000 508.470 504.000 ;
        RECT 508.230 499.450 508.370 500.000 ;
        RECT 508.170 499.130 508.430 499.450 ;
        RECT 508.400 498.110 508.660 498.430 ;
        RECT 508.460 492.650 508.600 498.110 ;
        RECT 508.400 492.330 508.660 492.650 ;
        RECT 530.940 491.650 531.200 491.970 ;
        RECT 531.000 487.890 531.140 491.650 ;
        RECT 530.940 487.570 531.200 487.890 ;
        RECT 570.500 487.570 570.760 487.890 ;
        RECT 570.560 182.230 570.700 487.570 ;
        RECT 570.500 181.910 570.760 182.230 ;
        RECT 924.700 181.910 924.960 182.230 ;
        RECT 924.760 2.400 924.900 181.910 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.570 500.000 509.850 504.000 ;
        RECT 509.610 498.680 509.750 500.000 ;
        RECT 509.380 498.540 509.750 498.680 ;
        RECT 509.380 484.005 509.520 498.540 ;
        RECT 509.310 483.635 509.590 484.005 ;
        RECT 938.490 101.475 938.770 101.845 ;
        RECT 938.560 82.870 938.700 101.475 ;
        RECT 938.560 82.730 942.840 82.870 ;
        RECT 942.700 2.400 942.840 82.730 ;
        RECT 942.490 -4.800 943.050 2.400 ;
      LAYER via2 ;
        RECT 509.310 483.680 509.590 483.960 ;
        RECT 938.490 101.520 938.770 101.800 ;
      LAYER met3 ;
        RECT 509.285 483.980 509.615 483.985 ;
        RECT 509.030 483.970 509.615 483.980 ;
        RECT 508.830 483.670 509.615 483.970 ;
        RECT 509.030 483.660 509.615 483.670 ;
        RECT 509.285 483.655 509.615 483.660 ;
        RECT 509.030 101.810 509.410 101.820 ;
        RECT 938.465 101.810 938.795 101.825 ;
        RECT 509.030 101.510 938.795 101.810 ;
        RECT 509.030 101.500 509.410 101.510 ;
        RECT 938.465 101.495 938.795 101.510 ;
      LAYER via3 ;
        RECT 509.060 483.660 509.380 483.980 ;
        RECT 509.060 101.500 509.380 101.820 ;
      LAYER met4 ;
        RECT 509.055 483.655 509.385 483.985 ;
        RECT 509.070 101.825 509.370 483.655 ;
        RECT 509.055 101.495 509.385 101.825 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 509.750 496.640 510.070 496.700 ;
        RECT 515.270 496.640 515.590 496.700 ;
        RECT 509.750 496.500 515.590 496.640 ;
        RECT 509.750 496.440 510.070 496.500 ;
        RECT 515.270 496.440 515.590 496.500 ;
        RECT 513.430 464.680 513.750 464.740 ;
        RECT 515.270 464.680 515.590 464.740 ;
        RECT 513.430 464.540 515.590 464.680 ;
        RECT 513.430 464.480 513.750 464.540 ;
        RECT 515.270 464.480 515.590 464.540 ;
        RECT 513.430 144.060 513.750 144.120 ;
        RECT 959.170 144.060 959.490 144.120 ;
        RECT 513.430 143.920 959.490 144.060 ;
        RECT 513.430 143.860 513.750 143.920 ;
        RECT 959.170 143.860 959.490 143.920 ;
      LAYER via ;
        RECT 509.780 496.440 510.040 496.700 ;
        RECT 515.300 496.440 515.560 496.700 ;
        RECT 513.460 464.480 513.720 464.740 ;
        RECT 515.300 464.480 515.560 464.740 ;
        RECT 513.460 143.860 513.720 144.120 ;
        RECT 959.200 143.860 959.460 144.120 ;
      LAYER met2 ;
        RECT 510.950 500.000 511.230 504.000 ;
        RECT 510.990 498.680 511.130 500.000 ;
        RECT 510.760 498.540 511.130 498.680 ;
        RECT 510.760 498.170 510.900 498.540 ;
        RECT 509.840 498.030 510.900 498.170 ;
        RECT 509.840 496.730 509.980 498.030 ;
        RECT 509.780 496.410 510.040 496.730 ;
        RECT 515.300 496.410 515.560 496.730 ;
        RECT 515.360 464.770 515.500 496.410 ;
        RECT 513.460 464.450 513.720 464.770 ;
        RECT 515.300 464.450 515.560 464.770 ;
        RECT 513.520 144.150 513.660 464.450 ;
        RECT 513.460 143.830 513.720 144.150 ;
        RECT 959.200 143.830 959.460 144.150 ;
        RECT 959.260 82.870 959.400 143.830 ;
        RECT 959.260 82.730 960.320 82.870 ;
        RECT 960.180 2.400 960.320 82.730 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.590 473.180 511.910 473.240 ;
        RECT 514.350 473.180 514.670 473.240 ;
        RECT 511.590 473.040 514.670 473.180 ;
        RECT 511.590 472.980 511.910 473.040 ;
        RECT 514.350 472.980 514.670 473.040 ;
        RECT 514.350 186.220 514.670 186.280 ;
        RECT 972.970 186.220 973.290 186.280 ;
        RECT 514.350 186.080 973.290 186.220 ;
        RECT 514.350 186.020 514.670 186.080 ;
        RECT 972.970 186.020 973.290 186.080 ;
      LAYER via ;
        RECT 511.620 472.980 511.880 473.240 ;
        RECT 514.380 472.980 514.640 473.240 ;
        RECT 514.380 186.020 514.640 186.280 ;
        RECT 973.000 186.020 973.260 186.280 ;
      LAYER met2 ;
        RECT 512.330 500.000 512.610 504.000 ;
        RECT 512.370 498.850 512.510 500.000 ;
        RECT 512.140 498.710 512.510 498.850 ;
        RECT 512.140 498.680 512.280 498.710 ;
        RECT 511.680 498.540 512.280 498.680 ;
        RECT 511.680 473.270 511.820 498.540 ;
        RECT 511.620 472.950 511.880 473.270 ;
        RECT 514.380 472.950 514.640 473.270 ;
        RECT 514.440 186.310 514.580 472.950 ;
        RECT 514.380 185.990 514.640 186.310 ;
        RECT 973.000 185.990 973.260 186.310 ;
        RECT 973.060 82.870 973.200 185.990 ;
        RECT 973.060 82.730 975.960 82.870 ;
        RECT 975.820 1.770 975.960 82.730 ;
        RECT 977.910 1.770 978.470 2.400 ;
        RECT 975.820 1.630 978.470 1.770 ;
        RECT 977.910 -4.800 978.470 1.630 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 487.440 499.500 487.760 499.760 ;
        RECT 487.530 497.720 487.670 499.500 ;
        RECT 487.210 497.520 487.670 497.720 ;
        RECT 487.210 497.460 487.530 497.520 ;
        RECT 485.370 473.520 485.690 473.580 ;
        RECT 487.210 473.520 487.530 473.580 ;
        RECT 485.370 473.380 487.530 473.520 ;
        RECT 485.370 473.320 485.690 473.380 ;
        RECT 487.210 473.320 487.530 473.380 ;
        RECT 485.370 24.720 485.690 24.780 ;
        RECT 658.790 24.720 659.110 24.780 ;
        RECT 485.370 24.580 659.110 24.720 ;
        RECT 485.370 24.520 485.690 24.580 ;
        RECT 658.790 24.520 659.110 24.580 ;
      LAYER via ;
        RECT 487.470 499.500 487.730 499.760 ;
        RECT 487.240 497.460 487.500 497.720 ;
        RECT 485.400 473.320 485.660 473.580 ;
        RECT 487.240 473.320 487.500 473.580 ;
        RECT 485.400 24.520 485.660 24.780 ;
        RECT 658.820 24.520 659.080 24.780 ;
      LAYER met2 ;
        RECT 487.490 500.000 487.770 504.000 ;
        RECT 487.530 499.790 487.670 500.000 ;
        RECT 487.470 499.470 487.730 499.790 ;
        RECT 487.240 497.430 487.500 497.750 ;
        RECT 487.300 473.610 487.440 497.430 ;
        RECT 485.400 473.290 485.660 473.610 ;
        RECT 487.240 473.290 487.500 473.610 ;
        RECT 485.460 24.810 485.600 473.290 ;
        RECT 485.400 24.490 485.660 24.810 ;
        RECT 658.820 24.490 659.080 24.810 ;
        RECT 658.880 2.400 659.020 24.490 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 513.890 164.460 514.210 164.520 ;
        RECT 993.670 164.460 993.990 164.520 ;
        RECT 513.890 164.320 993.990 164.460 ;
        RECT 513.890 164.260 514.210 164.320 ;
        RECT 993.670 164.260 993.990 164.320 ;
      LAYER via ;
        RECT 513.920 164.260 514.180 164.520 ;
        RECT 993.700 164.260 993.960 164.520 ;
      LAYER met2 ;
        RECT 513.710 500.000 513.990 504.000 ;
        RECT 513.750 498.850 513.890 500.000 ;
        RECT 513.750 498.710 514.120 498.850 ;
        RECT 513.980 164.550 514.120 498.710 ;
        RECT 513.920 164.230 514.180 164.550 ;
        RECT 993.700 164.230 993.960 164.550 ;
        RECT 993.760 1.770 993.900 164.230 ;
        RECT 995.390 1.770 995.950 2.400 ;
        RECT 993.760 1.630 995.950 1.770 ;
        RECT 995.390 -4.800 995.950 1.630 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1007.470 58.380 1007.790 58.440 ;
        RECT 1013.450 58.380 1013.770 58.440 ;
        RECT 1007.470 58.240 1013.770 58.380 ;
        RECT 1007.470 58.180 1007.790 58.240 ;
        RECT 1013.450 58.180 1013.770 58.240 ;
      LAYER via ;
        RECT 1007.500 58.180 1007.760 58.440 ;
        RECT 1013.480 58.180 1013.740 58.440 ;
      LAYER met2 ;
        RECT 515.090 500.000 515.370 504.000 ;
        RECT 515.130 498.340 515.270 500.000 ;
        RECT 514.900 498.200 515.270 498.340 ;
        RECT 514.900 484.005 515.040 498.200 ;
        RECT 514.830 483.635 515.110 484.005 ;
        RECT 1007.490 148.395 1007.770 148.765 ;
        RECT 1007.560 58.470 1007.700 148.395 ;
        RECT 1007.500 58.150 1007.760 58.470 ;
        RECT 1013.480 58.150 1013.740 58.470 ;
        RECT 1013.540 2.400 1013.680 58.150 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
      LAYER via2 ;
        RECT 514.830 483.680 515.110 483.960 ;
        RECT 1007.490 148.440 1007.770 148.720 ;
      LAYER met3 ;
        RECT 513.630 483.970 514.010 483.980 ;
        RECT 514.805 483.970 515.135 483.985 ;
        RECT 513.630 483.670 515.135 483.970 ;
        RECT 513.630 483.660 514.010 483.670 ;
        RECT 514.805 483.655 515.135 483.670 ;
        RECT 513.630 148.730 514.010 148.740 ;
        RECT 1007.465 148.730 1007.795 148.745 ;
        RECT 513.630 148.430 1007.795 148.730 ;
        RECT 513.630 148.420 514.010 148.430 ;
        RECT 1007.465 148.415 1007.795 148.430 ;
      LAYER via3 ;
        RECT 513.660 483.660 513.980 483.980 ;
        RECT 513.660 148.420 513.980 148.740 ;
      LAYER met4 ;
        RECT 513.655 483.655 513.985 483.985 ;
        RECT 513.670 148.745 513.970 483.655 ;
        RECT 513.655 148.415 513.985 148.745 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 516.420 498.820 516.740 499.080 ;
        RECT 516.510 498.400 516.650 498.820 ;
        RECT 516.510 498.200 516.970 498.400 ;
        RECT 516.650 498.140 516.970 498.200 ;
        RECT 516.650 486.100 516.970 486.160 ;
        RECT 578.750 486.100 579.070 486.160 ;
        RECT 516.650 485.960 579.070 486.100 ;
        RECT 516.650 485.900 516.970 485.960 ;
        RECT 578.750 485.900 579.070 485.960 ;
        RECT 577.830 182.480 578.150 182.540 ;
        RECT 1028.170 182.480 1028.490 182.540 ;
        RECT 577.830 182.340 1028.490 182.480 ;
        RECT 577.830 182.280 578.150 182.340 ;
        RECT 1028.170 182.280 1028.490 182.340 ;
      LAYER via ;
        RECT 516.450 498.820 516.710 499.080 ;
        RECT 516.680 498.140 516.940 498.400 ;
        RECT 516.680 485.900 516.940 486.160 ;
        RECT 578.780 485.900 579.040 486.160 ;
        RECT 577.860 182.280 578.120 182.540 ;
        RECT 1028.200 182.280 1028.460 182.540 ;
      LAYER met2 ;
        RECT 516.470 500.000 516.750 504.000 ;
        RECT 516.510 499.110 516.650 500.000 ;
        RECT 516.450 498.790 516.710 499.110 ;
        RECT 516.680 498.110 516.940 498.430 ;
        RECT 516.740 486.190 516.880 498.110 ;
        RECT 516.680 485.870 516.940 486.190 ;
        RECT 578.780 485.870 579.040 486.190 ;
        RECT 578.840 420.970 578.980 485.870 ;
        RECT 577.920 420.830 578.980 420.970 ;
        RECT 577.920 182.570 578.060 420.830 ;
        RECT 577.860 182.250 578.120 182.570 ;
        RECT 1028.200 182.250 1028.460 182.570 ;
        RECT 1028.260 82.870 1028.400 182.250 ;
        RECT 1028.260 82.730 1031.160 82.870 ;
        RECT 1031.020 2.400 1031.160 82.730 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.800 499.500 518.120 499.760 ;
        RECT 517.890 496.640 518.030 499.500 ;
        RECT 522.630 496.640 522.950 496.700 ;
        RECT 517.890 496.500 522.950 496.640 ;
        RECT 522.630 496.440 522.950 496.500 ;
        RECT 521.710 185.880 522.030 185.940 ;
        RECT 1049.330 185.880 1049.650 185.940 ;
        RECT 521.710 185.740 1049.650 185.880 ;
        RECT 521.710 185.680 522.030 185.740 ;
        RECT 1049.330 185.680 1049.650 185.740 ;
      LAYER via ;
        RECT 517.830 499.500 518.090 499.760 ;
        RECT 522.660 496.440 522.920 496.700 ;
        RECT 521.740 185.680 522.000 185.940 ;
        RECT 1049.360 185.680 1049.620 185.940 ;
      LAYER met2 ;
        RECT 517.850 500.000 518.130 504.000 ;
        RECT 517.890 499.790 518.030 500.000 ;
        RECT 517.830 499.470 518.090 499.790 ;
        RECT 522.660 496.410 522.920 496.730 ;
        RECT 522.720 420.970 522.860 496.410 ;
        RECT 521.800 420.830 522.860 420.970 ;
        RECT 521.800 185.970 521.940 420.830 ;
        RECT 521.740 185.650 522.000 185.970 ;
        RECT 1049.360 185.650 1049.620 185.970 ;
        RECT 1049.420 34.570 1049.560 185.650 ;
        RECT 1048.960 34.430 1049.560 34.570 ;
        RECT 1048.960 2.400 1049.100 34.430 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 519.180 499.500 519.500 499.760 ;
        RECT 519.270 497.320 519.410 499.500 ;
        RECT 520.330 497.320 520.650 497.380 ;
        RECT 519.270 497.180 520.650 497.320 ;
        RECT 520.330 497.120 520.650 497.180 ;
        RECT 520.330 151.200 520.650 151.260 ;
        RECT 1062.670 151.200 1062.990 151.260 ;
        RECT 520.330 151.060 1062.990 151.200 ;
        RECT 520.330 151.000 520.650 151.060 ;
        RECT 1062.670 151.000 1062.990 151.060 ;
      LAYER via ;
        RECT 519.210 499.500 519.470 499.760 ;
        RECT 520.360 497.120 520.620 497.380 ;
        RECT 520.360 151.000 520.620 151.260 ;
        RECT 1062.700 151.000 1062.960 151.260 ;
      LAYER met2 ;
        RECT 519.230 500.000 519.510 504.000 ;
        RECT 519.270 499.790 519.410 500.000 ;
        RECT 519.210 499.470 519.470 499.790 ;
        RECT 520.360 497.090 520.620 497.410 ;
        RECT 520.420 151.290 520.560 497.090 ;
        RECT 520.360 150.970 520.620 151.290 ;
        RECT 1062.700 150.970 1062.960 151.290 ;
        RECT 1062.760 82.870 1062.900 150.970 ;
        RECT 1062.760 82.730 1067.040 82.870 ;
        RECT 1066.900 2.400 1067.040 82.730 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 520.790 150.860 521.110 150.920 ;
        RECT 1083.370 150.860 1083.690 150.920 ;
        RECT 520.790 150.720 1083.690 150.860 ;
        RECT 520.790 150.660 521.110 150.720 ;
        RECT 1083.370 150.660 1083.690 150.720 ;
      LAYER via ;
        RECT 520.820 150.660 521.080 150.920 ;
        RECT 1083.400 150.660 1083.660 150.920 ;
      LAYER met2 ;
        RECT 520.610 500.000 520.890 504.000 ;
        RECT 520.650 498.340 520.790 500.000 ;
        RECT 520.650 498.200 521.020 498.340 ;
        RECT 520.880 150.950 521.020 498.200 ;
        RECT 520.820 150.630 521.080 150.950 ;
        RECT 1083.400 150.630 1083.660 150.950 ;
        RECT 1083.460 82.870 1083.600 150.630 ;
        RECT 1083.460 82.730 1084.520 82.870 ;
        RECT 1084.380 2.400 1084.520 82.730 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 521.940 498.820 522.260 499.080 ;
        RECT 522.030 497.720 522.170 498.820 ;
        RECT 521.710 497.520 522.170 497.720 ;
        RECT 521.710 497.460 522.030 497.520 ;
        RECT 521.250 164.120 521.570 164.180 ;
        RECT 1097.170 164.120 1097.490 164.180 ;
        RECT 521.250 163.980 1097.490 164.120 ;
        RECT 521.250 163.920 521.570 163.980 ;
        RECT 1097.170 163.920 1097.490 163.980 ;
      LAYER via ;
        RECT 521.970 498.820 522.230 499.080 ;
        RECT 521.740 497.460 522.000 497.720 ;
        RECT 521.280 163.920 521.540 164.180 ;
        RECT 1097.200 163.920 1097.460 164.180 ;
      LAYER met2 ;
        RECT 521.990 500.000 522.270 504.000 ;
        RECT 522.030 499.110 522.170 500.000 ;
        RECT 521.970 498.790 522.230 499.110 ;
        RECT 521.740 497.430 522.000 497.750 ;
        RECT 521.800 476.170 521.940 497.430 ;
        RECT 521.340 476.030 521.940 476.170 ;
        RECT 521.340 164.210 521.480 476.030 ;
        RECT 521.280 163.890 521.540 164.210 ;
        RECT 1097.200 163.890 1097.460 164.210 ;
        RECT 1097.260 82.870 1097.400 163.890 ;
        RECT 1097.260 82.730 1100.160 82.870 ;
        RECT 1100.020 1.770 1100.160 82.730 ;
        RECT 1102.110 1.770 1102.670 2.400 ;
        RECT 1100.020 1.630 1102.670 1.770 ;
        RECT 1102.110 -4.800 1102.670 1.630 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.370 500.000 523.650 504.000 ;
        RECT 523.410 498.850 523.550 500.000 ;
        RECT 523.410 498.710 523.780 498.850 ;
        RECT 523.640 486.045 523.780 498.710 ;
        RECT 523.570 485.675 523.850 486.045 ;
        RECT 1117.890 147.715 1118.170 148.085 ;
        RECT 1117.960 1.770 1118.100 147.715 ;
        RECT 1119.590 1.770 1120.150 2.400 ;
        RECT 1117.960 1.630 1120.150 1.770 ;
        RECT 1119.590 -4.800 1120.150 1.630 ;
      LAYER via2 ;
        RECT 523.570 485.720 523.850 486.000 ;
        RECT 1117.890 147.760 1118.170 148.040 ;
      LAYER met3 ;
        RECT 520.990 486.010 521.370 486.020 ;
        RECT 523.545 486.010 523.875 486.025 ;
        RECT 520.990 485.710 523.875 486.010 ;
        RECT 520.990 485.700 521.370 485.710 ;
        RECT 523.545 485.695 523.875 485.710 ;
        RECT 520.990 148.050 521.370 148.060 ;
        RECT 1117.865 148.050 1118.195 148.065 ;
        RECT 520.990 147.750 1118.195 148.050 ;
        RECT 520.990 147.740 521.370 147.750 ;
        RECT 1117.865 147.735 1118.195 147.750 ;
      LAYER via3 ;
        RECT 521.020 485.700 521.340 486.020 ;
        RECT 521.020 147.740 521.340 148.060 ;
      LAYER met4 ;
        RECT 521.015 485.695 521.345 486.025 ;
        RECT 521.030 148.065 521.330 485.695 ;
        RECT 521.015 147.735 521.345 148.065 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.700 499.500 525.020 499.760 ;
        RECT 524.790 497.320 524.930 499.500 ;
        RECT 529.070 497.320 529.390 497.380 ;
        RECT 524.790 497.180 529.390 497.320 ;
        RECT 529.070 497.120 529.390 497.180 ;
        RECT 528.610 171.600 528.930 171.660 ;
        RECT 1131.670 171.600 1131.990 171.660 ;
        RECT 528.610 171.460 1131.990 171.600 ;
        RECT 528.610 171.400 528.930 171.460 ;
        RECT 1131.670 171.400 1131.990 171.460 ;
        RECT 1131.670 19.280 1131.990 19.340 ;
        RECT 1137.650 19.280 1137.970 19.340 ;
        RECT 1131.670 19.140 1137.970 19.280 ;
        RECT 1131.670 19.080 1131.990 19.140 ;
        RECT 1137.650 19.080 1137.970 19.140 ;
      LAYER via ;
        RECT 524.730 499.500 524.990 499.760 ;
        RECT 529.100 497.120 529.360 497.380 ;
        RECT 528.640 171.400 528.900 171.660 ;
        RECT 1131.700 171.400 1131.960 171.660 ;
        RECT 1131.700 19.080 1131.960 19.340 ;
        RECT 1137.680 19.080 1137.940 19.340 ;
      LAYER met2 ;
        RECT 524.750 500.000 525.030 504.000 ;
        RECT 524.790 499.790 524.930 500.000 ;
        RECT 524.730 499.470 524.990 499.790 ;
        RECT 529.100 497.090 529.360 497.410 ;
        RECT 529.160 420.970 529.300 497.090 ;
        RECT 528.700 420.830 529.300 420.970 ;
        RECT 528.700 171.690 528.840 420.830 ;
        RECT 528.640 171.370 528.900 171.690 ;
        RECT 1131.700 171.370 1131.960 171.690 ;
        RECT 1131.760 19.370 1131.900 171.370 ;
        RECT 1131.700 19.050 1131.960 19.370 ;
        RECT 1137.680 19.050 1137.940 19.370 ;
        RECT 1137.740 2.400 1137.880 19.050 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 526.080 499.500 526.400 499.760 ;
        RECT 526.170 498.060 526.310 499.500 ;
        RECT 525.850 497.860 526.310 498.060 ;
        RECT 525.850 497.800 526.170 497.860 ;
        RECT 525.850 488.140 526.170 488.200 ;
        RECT 527.230 488.140 527.550 488.200 ;
        RECT 525.850 488.000 527.550 488.140 ;
        RECT 525.850 487.940 526.170 488.000 ;
        RECT 527.230 487.940 527.550 488.000 ;
        RECT 527.230 154.600 527.550 154.660 ;
        RECT 1152.370 154.600 1152.690 154.660 ;
        RECT 527.230 154.460 1152.690 154.600 ;
        RECT 527.230 154.400 527.550 154.460 ;
        RECT 1152.370 154.400 1152.690 154.460 ;
      LAYER via ;
        RECT 526.110 499.500 526.370 499.760 ;
        RECT 525.880 497.800 526.140 498.060 ;
        RECT 525.880 487.940 526.140 488.200 ;
        RECT 527.260 487.940 527.520 488.200 ;
        RECT 527.260 154.400 527.520 154.660 ;
        RECT 1152.400 154.400 1152.660 154.660 ;
      LAYER met2 ;
        RECT 526.130 500.000 526.410 504.000 ;
        RECT 526.170 499.790 526.310 500.000 ;
        RECT 526.110 499.470 526.370 499.790 ;
        RECT 525.880 497.770 526.140 498.090 ;
        RECT 525.940 488.230 526.080 497.770 ;
        RECT 525.880 487.910 526.140 488.230 ;
        RECT 527.260 487.910 527.520 488.230 ;
        RECT 527.320 154.690 527.460 487.910 ;
        RECT 527.260 154.370 527.520 154.690 ;
        RECT 1152.400 154.370 1152.660 154.690 ;
        RECT 1152.460 82.870 1152.600 154.370 ;
        RECT 1152.460 82.730 1155.360 82.870 ;
        RECT 1155.220 2.400 1155.360 82.730 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 488.820 499.500 489.140 499.760 ;
        RECT 488.910 498.740 489.050 499.500 ;
        RECT 488.590 498.540 489.050 498.740 ;
        RECT 488.590 498.480 488.910 498.540 ;
      LAYER via ;
        RECT 488.850 499.500 489.110 499.760 ;
        RECT 488.620 498.480 488.880 498.740 ;
      LAYER met2 ;
        RECT 488.870 500.000 489.150 504.000 ;
        RECT 488.910 499.790 489.050 500.000 ;
        RECT 488.850 499.470 489.110 499.790 ;
        RECT 488.620 498.450 488.880 498.770 ;
        RECT 488.680 498.285 488.820 498.450 ;
        RECT 488.610 497.915 488.890 498.285 ;
        RECT 676.750 122.555 677.030 122.925 ;
        RECT 676.820 34.570 676.960 122.555 ;
        RECT 676.360 34.430 676.960 34.570 ;
        RECT 676.360 2.400 676.500 34.430 ;
        RECT 676.150 -4.800 676.710 2.400 ;
      LAYER via2 ;
        RECT 488.610 497.960 488.890 498.240 ;
        RECT 676.750 122.600 677.030 122.880 ;
      LAYER met3 ;
        RECT 486.950 498.250 487.330 498.260 ;
        RECT 488.585 498.250 488.915 498.265 ;
        RECT 486.950 497.950 488.915 498.250 ;
        RECT 486.950 497.940 487.330 497.950 ;
        RECT 488.585 497.935 488.915 497.950 ;
        RECT 486.950 122.890 487.330 122.900 ;
        RECT 676.725 122.890 677.055 122.905 ;
        RECT 486.950 122.590 677.055 122.890 ;
        RECT 486.950 122.580 487.330 122.590 ;
        RECT 676.725 122.575 677.055 122.590 ;
      LAYER via3 ;
        RECT 486.980 497.940 487.300 498.260 ;
        RECT 486.980 122.580 487.300 122.900 ;
      LAYER met4 ;
        RECT 486.975 497.935 487.305 498.265 ;
        RECT 486.990 122.905 487.290 497.935 ;
        RECT 486.975 122.575 487.305 122.905 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.460 499.500 527.780 499.760 ;
        RECT 527.550 498.340 527.690 499.500 ;
        RECT 528.150 498.340 528.470 498.400 ;
        RECT 527.550 498.200 528.470 498.340 ;
        RECT 528.150 498.140 528.470 498.200 ;
        RECT 528.150 154.940 528.470 155.000 ;
        RECT 1173.070 154.940 1173.390 155.000 ;
        RECT 528.150 154.800 1173.390 154.940 ;
        RECT 528.150 154.740 528.470 154.800 ;
        RECT 1173.070 154.740 1173.390 154.800 ;
      LAYER via ;
        RECT 527.490 499.500 527.750 499.760 ;
        RECT 528.180 498.140 528.440 498.400 ;
        RECT 528.180 154.740 528.440 155.000 ;
        RECT 1173.100 154.740 1173.360 155.000 ;
      LAYER met2 ;
        RECT 527.510 500.000 527.790 504.000 ;
        RECT 527.550 499.790 527.690 500.000 ;
        RECT 527.490 499.470 527.750 499.790 ;
        RECT 528.180 498.110 528.440 498.430 ;
        RECT 528.240 155.030 528.380 498.110 ;
        RECT 528.180 154.710 528.440 155.030 ;
        RECT 1173.100 154.710 1173.360 155.030 ;
        RECT 1173.160 2.400 1173.300 154.710 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 528.840 499.500 529.160 499.760 ;
        RECT 528.930 499.020 529.070 499.500 ;
        RECT 528.930 498.880 529.300 499.020 ;
        RECT 529.160 498.400 529.300 498.880 ;
        RECT 529.070 498.140 529.390 498.400 ;
        RECT 527.690 472.840 528.010 472.900 ;
        RECT 528.610 472.840 528.930 472.900 ;
        RECT 527.690 472.700 528.930 472.840 ;
        RECT 527.690 472.640 528.010 472.700 ;
        RECT 528.610 472.640 528.930 472.700 ;
        RECT 527.690 158.680 528.010 158.740 ;
        RECT 1186.870 158.680 1187.190 158.740 ;
        RECT 527.690 158.540 1187.190 158.680 ;
        RECT 527.690 158.480 528.010 158.540 ;
        RECT 1186.870 158.480 1187.190 158.540 ;
      LAYER via ;
        RECT 528.870 499.500 529.130 499.760 ;
        RECT 529.100 498.140 529.360 498.400 ;
        RECT 527.720 472.640 527.980 472.900 ;
        RECT 528.640 472.640 528.900 472.900 ;
        RECT 527.720 158.480 527.980 158.740 ;
        RECT 1186.900 158.480 1187.160 158.740 ;
      LAYER met2 ;
        RECT 528.890 500.000 529.170 504.000 ;
        RECT 528.930 499.790 529.070 500.000 ;
        RECT 528.870 499.470 529.130 499.790 ;
        RECT 529.100 498.340 529.360 498.430 ;
        RECT 528.700 498.200 529.360 498.340 ;
        RECT 528.700 472.930 528.840 498.200 ;
        RECT 529.100 498.110 529.360 498.200 ;
        RECT 527.720 472.610 527.980 472.930 ;
        RECT 528.640 472.610 528.900 472.930 ;
        RECT 527.780 158.770 527.920 472.610 ;
        RECT 527.720 158.450 527.980 158.770 ;
        RECT 1186.900 158.450 1187.160 158.770 ;
        RECT 1186.960 82.870 1187.100 158.450 ;
        RECT 1186.960 82.730 1188.480 82.870 ;
        RECT 1188.340 1.770 1188.480 82.730 ;
        RECT 1190.430 1.770 1190.990 2.400 ;
        RECT 1188.340 1.630 1190.990 1.770 ;
        RECT 1190.430 -4.800 1190.990 1.630 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 530.220 499.700 530.540 499.760 ;
        RECT 530.080 499.500 530.540 499.700 ;
        RECT 530.080 499.080 530.220 499.500 ;
        RECT 529.990 498.820 530.310 499.080 ;
        RECT 529.990 485.420 530.310 485.480 ;
        RECT 584.270 485.420 584.590 485.480 ;
        RECT 529.990 485.280 584.590 485.420 ;
        RECT 529.990 485.220 530.310 485.280 ;
        RECT 584.270 485.220 584.590 485.280 ;
        RECT 584.730 185.540 585.050 185.600 ;
        RECT 1207.570 185.540 1207.890 185.600 ;
        RECT 584.730 185.400 1207.890 185.540 ;
        RECT 584.730 185.340 585.050 185.400 ;
        RECT 1207.570 185.340 1207.890 185.400 ;
      LAYER via ;
        RECT 530.250 499.500 530.510 499.760 ;
        RECT 530.020 498.820 530.280 499.080 ;
        RECT 530.020 485.220 530.280 485.480 ;
        RECT 584.300 485.220 584.560 485.480 ;
        RECT 584.760 185.340 585.020 185.600 ;
        RECT 1207.600 185.340 1207.860 185.600 ;
      LAYER met2 ;
        RECT 530.270 500.000 530.550 504.000 ;
        RECT 530.310 499.790 530.450 500.000 ;
        RECT 530.250 499.470 530.510 499.790 ;
        RECT 530.020 498.790 530.280 499.110 ;
        RECT 530.080 485.510 530.220 498.790 ;
        RECT 530.020 485.190 530.280 485.510 ;
        RECT 584.300 485.190 584.560 485.510 ;
        RECT 584.360 472.330 584.500 485.190 ;
        RECT 584.360 472.190 584.960 472.330 ;
        RECT 584.820 185.630 584.960 472.190 ;
        RECT 584.760 185.310 585.020 185.630 ;
        RECT 1207.600 185.310 1207.860 185.630 ;
        RECT 1207.660 82.870 1207.800 185.310 ;
        RECT 1207.660 82.730 1208.720 82.870 ;
        RECT 1208.580 2.400 1208.720 82.730 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.830 489.840 532.150 489.900 ;
        RECT 534.590 489.840 534.910 489.900 ;
        RECT 531.830 489.700 534.910 489.840 ;
        RECT 531.830 489.640 532.150 489.700 ;
        RECT 534.590 489.640 534.910 489.700 ;
        RECT 534.590 158.340 534.910 158.400 ;
        RECT 1221.370 158.340 1221.690 158.400 ;
        RECT 534.590 158.200 1221.690 158.340 ;
        RECT 534.590 158.140 534.910 158.200 ;
        RECT 1221.370 158.140 1221.690 158.200 ;
      LAYER via ;
        RECT 531.860 489.640 532.120 489.900 ;
        RECT 534.620 489.640 534.880 489.900 ;
        RECT 534.620 158.140 534.880 158.400 ;
        RECT 1221.400 158.140 1221.660 158.400 ;
      LAYER met2 ;
        RECT 531.650 500.000 531.930 504.000 ;
        RECT 531.690 498.340 531.830 500.000 ;
        RECT 531.690 498.200 532.060 498.340 ;
        RECT 531.920 489.930 532.060 498.200 ;
        RECT 531.860 489.610 532.120 489.930 ;
        RECT 534.620 489.610 534.880 489.930 ;
        RECT 534.680 158.430 534.820 489.610 ;
        RECT 534.620 158.110 534.880 158.430 ;
        RECT 1221.400 158.110 1221.660 158.430 ;
        RECT 1221.460 82.870 1221.600 158.110 ;
        RECT 1221.460 82.730 1226.200 82.870 ;
        RECT 1226.060 2.400 1226.200 82.730 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 535.510 184.860 535.830 184.920 ;
        RECT 1242.070 184.860 1242.390 184.920 ;
        RECT 535.510 184.720 1242.390 184.860 ;
        RECT 535.510 184.660 535.830 184.720 ;
        RECT 1242.070 184.660 1242.390 184.720 ;
      LAYER via ;
        RECT 535.540 184.660 535.800 184.920 ;
        RECT 1242.100 184.660 1242.360 184.920 ;
      LAYER met2 ;
        RECT 533.030 500.000 533.310 504.000 ;
        RECT 533.070 498.965 533.210 500.000 ;
        RECT 533.000 498.595 533.280 498.965 ;
        RECT 535.530 486.355 535.810 486.725 ;
        RECT 535.600 184.950 535.740 486.355 ;
        RECT 535.540 184.630 535.800 184.950 ;
        RECT 1242.100 184.630 1242.360 184.950 ;
        RECT 1242.160 1.770 1242.300 184.630 ;
        RECT 1243.790 1.770 1244.350 2.400 ;
        RECT 1242.160 1.630 1244.350 1.770 ;
        RECT 1243.790 -4.800 1244.350 1.630 ;
      LAYER via2 ;
        RECT 533.000 498.640 533.280 498.920 ;
        RECT 535.530 486.400 535.810 486.680 ;
      LAYER met3 ;
        RECT 532.975 498.940 533.305 498.945 ;
        RECT 532.950 498.930 533.330 498.940 ;
        RECT 532.520 498.630 533.330 498.930 ;
        RECT 532.950 498.620 533.330 498.630 ;
        RECT 532.975 498.615 533.305 498.620 ;
        RECT 532.950 486.690 533.330 486.700 ;
        RECT 535.505 486.690 535.835 486.705 ;
        RECT 532.950 486.390 535.835 486.690 ;
        RECT 532.950 486.380 533.330 486.390 ;
        RECT 535.505 486.375 535.835 486.390 ;
      LAYER via3 ;
        RECT 532.980 498.620 533.300 498.940 ;
        RECT 532.980 486.380 533.300 486.700 ;
      LAYER met4 ;
        RECT 532.975 498.615 533.305 498.945 ;
        RECT 532.990 486.705 533.290 498.615 ;
        RECT 532.975 486.375 533.305 486.705 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 534.360 499.500 534.680 499.760 ;
        RECT 533.210 498.000 533.530 498.060 ;
        RECT 534.450 498.000 534.590 499.500 ;
        RECT 533.210 497.860 534.590 498.000 ;
        RECT 533.210 497.800 533.530 497.860 ;
        RECT 533.210 488.140 533.530 488.200 ;
        RECT 535.050 488.140 535.370 488.200 ;
        RECT 533.210 488.000 535.370 488.140 ;
        RECT 533.210 487.940 533.530 488.000 ;
        RECT 535.050 487.940 535.370 488.000 ;
        RECT 535.050 158.000 535.370 158.060 ;
        RECT 1255.870 158.000 1256.190 158.060 ;
        RECT 535.050 157.860 1256.190 158.000 ;
        RECT 535.050 157.800 535.370 157.860 ;
        RECT 1255.870 157.800 1256.190 157.860 ;
        RECT 1255.870 18.940 1256.190 19.000 ;
        RECT 1261.850 18.940 1262.170 19.000 ;
        RECT 1255.870 18.800 1262.170 18.940 ;
        RECT 1255.870 18.740 1256.190 18.800 ;
        RECT 1261.850 18.740 1262.170 18.800 ;
      LAYER via ;
        RECT 534.390 499.500 534.650 499.760 ;
        RECT 533.240 497.800 533.500 498.060 ;
        RECT 533.240 487.940 533.500 488.200 ;
        RECT 535.080 487.940 535.340 488.200 ;
        RECT 535.080 157.800 535.340 158.060 ;
        RECT 1255.900 157.800 1256.160 158.060 ;
        RECT 1255.900 18.740 1256.160 19.000 ;
        RECT 1261.880 18.740 1262.140 19.000 ;
      LAYER met2 ;
        RECT 534.410 500.000 534.690 504.000 ;
        RECT 534.450 499.790 534.590 500.000 ;
        RECT 534.390 499.470 534.650 499.790 ;
        RECT 533.240 497.770 533.500 498.090 ;
        RECT 533.300 488.230 533.440 497.770 ;
        RECT 533.240 487.910 533.500 488.230 ;
        RECT 535.080 487.910 535.340 488.230 ;
        RECT 535.140 158.090 535.280 487.910 ;
        RECT 535.080 157.770 535.340 158.090 ;
        RECT 1255.900 157.770 1256.160 158.090 ;
        RECT 1255.960 19.030 1256.100 157.770 ;
        RECT 1255.900 18.710 1256.160 19.030 ;
        RECT 1261.880 18.710 1262.140 19.030 ;
        RECT 1261.940 2.400 1262.080 18.710 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 535.050 488.820 535.370 488.880 ;
        RECT 556.670 488.820 556.990 488.880 ;
        RECT 535.050 488.680 556.990 488.820 ;
        RECT 535.050 488.620 535.370 488.680 ;
        RECT 556.670 488.620 556.990 488.680 ;
        RECT 556.670 488.140 556.990 488.200 ;
        RECT 580.590 488.140 580.910 488.200 ;
        RECT 556.670 488.000 580.910 488.140 ;
        RECT 556.670 487.940 556.990 488.000 ;
        RECT 580.590 487.940 580.910 488.000 ;
        RECT 580.590 484.060 580.910 484.120 ;
        RECT 585.190 484.060 585.510 484.120 ;
        RECT 580.590 483.920 585.510 484.060 ;
        RECT 580.590 483.860 580.910 483.920 ;
        RECT 585.190 483.860 585.510 483.920 ;
        RECT 584.270 471.820 584.590 471.880 ;
        RECT 585.190 471.820 585.510 471.880 ;
        RECT 584.270 471.680 585.510 471.820 ;
        RECT 584.270 471.620 584.590 471.680 ;
        RECT 585.190 471.620 585.510 471.680 ;
        RECT 584.270 185.200 584.590 185.260 ;
        RECT 1276.570 185.200 1276.890 185.260 ;
        RECT 584.270 185.060 1276.890 185.200 ;
        RECT 584.270 185.000 584.590 185.060 ;
        RECT 1276.570 185.000 1276.890 185.060 ;
      LAYER via ;
        RECT 535.080 488.620 535.340 488.880 ;
        RECT 556.700 488.620 556.960 488.880 ;
        RECT 556.700 487.940 556.960 488.200 ;
        RECT 580.620 487.940 580.880 488.200 ;
        RECT 580.620 483.860 580.880 484.120 ;
        RECT 585.220 483.860 585.480 484.120 ;
        RECT 584.300 471.620 584.560 471.880 ;
        RECT 585.220 471.620 585.480 471.880 ;
        RECT 584.300 185.000 584.560 185.260 ;
        RECT 1276.600 185.000 1276.860 185.260 ;
      LAYER met2 ;
        RECT 535.790 500.000 536.070 504.000 ;
        RECT 535.830 499.020 535.970 500.000 ;
        RECT 535.140 498.880 535.970 499.020 ;
        RECT 535.140 488.910 535.280 498.880 ;
        RECT 535.080 488.590 535.340 488.910 ;
        RECT 556.700 488.590 556.960 488.910 ;
        RECT 556.760 488.230 556.900 488.590 ;
        RECT 556.700 487.910 556.960 488.230 ;
        RECT 580.620 487.910 580.880 488.230 ;
        RECT 580.680 484.150 580.820 487.910 ;
        RECT 580.620 483.830 580.880 484.150 ;
        RECT 585.220 483.830 585.480 484.150 ;
        RECT 585.280 471.910 585.420 483.830 ;
        RECT 584.300 471.590 584.560 471.910 ;
        RECT 585.220 471.590 585.480 471.910 ;
        RECT 584.360 185.290 584.500 471.590 ;
        RECT 584.300 184.970 584.560 185.290 ;
        RECT 1276.600 184.970 1276.860 185.290 ;
        RECT 1276.660 82.870 1276.800 184.970 ;
        RECT 1276.660 82.730 1279.560 82.870 ;
        RECT 1279.420 2.400 1279.560 82.730 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.170 500.000 537.450 504.000 ;
        RECT 537.210 499.815 537.350 500.000 ;
        RECT 537.140 499.445 537.420 499.815 ;
        RECT 1297.290 154.515 1297.570 154.885 ;
        RECT 1297.360 2.400 1297.500 154.515 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
      LAYER via2 ;
        RECT 537.140 499.490 537.420 499.770 ;
        RECT 1297.290 154.560 1297.570 154.840 ;
      LAYER met3 ;
        RECT 537.115 499.780 537.445 499.795 ;
        RECT 534.790 499.610 535.170 499.620 ;
        RECT 537.115 499.610 537.660 499.780 ;
        RECT 534.790 499.310 537.660 499.610 ;
        RECT 534.790 499.300 535.170 499.310 ;
        RECT 534.790 154.850 535.170 154.860 ;
        RECT 1297.265 154.850 1297.595 154.865 ;
        RECT 534.790 154.550 1297.595 154.850 ;
        RECT 534.790 154.540 535.170 154.550 ;
        RECT 1297.265 154.535 1297.595 154.550 ;
      LAYER via3 ;
        RECT 534.820 499.300 535.140 499.620 ;
        RECT 534.820 154.540 535.140 154.860 ;
      LAYER met4 ;
        RECT 534.815 499.295 535.145 499.625 ;
        RECT 534.830 154.865 535.130 499.295 ;
        RECT 534.815 154.535 535.145 154.865 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.500 499.500 538.820 499.760 ;
        RECT 538.590 498.740 538.730 499.500 ;
        RECT 538.590 498.540 539.050 498.740 ;
        RECT 538.730 498.480 539.050 498.540 ;
        RECT 539.190 472.980 539.510 473.240 ;
        RECT 539.280 471.140 539.420 472.980 ;
        RECT 539.280 471.000 541.720 471.140 ;
        RECT 541.580 470.860 541.720 471.000 ;
        RECT 541.490 470.600 541.810 470.860 ;
        RECT 541.490 184.520 541.810 184.580 ;
        RECT 1311.070 184.520 1311.390 184.580 ;
        RECT 541.490 184.380 1311.390 184.520 ;
        RECT 541.490 184.320 541.810 184.380 ;
        RECT 1311.070 184.320 1311.390 184.380 ;
      LAYER via ;
        RECT 538.530 499.500 538.790 499.760 ;
        RECT 538.760 498.480 539.020 498.740 ;
        RECT 539.220 472.980 539.480 473.240 ;
        RECT 541.520 470.600 541.780 470.860 ;
        RECT 541.520 184.320 541.780 184.580 ;
        RECT 1311.100 184.320 1311.360 184.580 ;
      LAYER met2 ;
        RECT 538.550 500.000 538.830 504.000 ;
        RECT 538.590 499.790 538.730 500.000 ;
        RECT 538.530 499.470 538.790 499.790 ;
        RECT 538.760 498.680 539.020 498.770 ;
        RECT 538.760 498.540 539.420 498.680 ;
        RECT 538.760 498.450 539.020 498.540 ;
        RECT 539.280 473.270 539.420 498.540 ;
        RECT 539.220 472.950 539.480 473.270 ;
        RECT 541.520 470.570 541.780 470.890 ;
        RECT 541.580 184.610 541.720 470.570 ;
        RECT 541.520 184.290 541.780 184.610 ;
        RECT 1311.100 184.290 1311.360 184.610 ;
        RECT 1311.160 82.870 1311.300 184.290 ;
        RECT 1311.160 82.730 1312.680 82.870 ;
        RECT 1312.540 1.770 1312.680 82.730 ;
        RECT 1314.630 1.770 1315.190 2.400 ;
        RECT 1312.540 1.630 1315.190 1.770 ;
        RECT 1314.630 -4.800 1315.190 1.630 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 539.650 491.540 539.970 491.600 ;
        RECT 541.030 491.540 541.350 491.600 ;
        RECT 539.650 491.400 541.350 491.540 ;
        RECT 539.650 491.340 539.970 491.400 ;
        RECT 541.030 491.340 541.350 491.400 ;
        RECT 541.030 163.780 541.350 163.840 ;
        RECT 1331.770 163.780 1332.090 163.840 ;
        RECT 541.030 163.640 1332.090 163.780 ;
        RECT 541.030 163.580 541.350 163.640 ;
        RECT 1331.770 163.580 1332.090 163.640 ;
      LAYER via ;
        RECT 539.680 491.340 539.940 491.600 ;
        RECT 541.060 491.340 541.320 491.600 ;
        RECT 541.060 163.580 541.320 163.840 ;
        RECT 1331.800 163.580 1332.060 163.840 ;
      LAYER met2 ;
        RECT 539.930 500.000 540.210 504.000 ;
        RECT 539.970 498.850 540.110 500.000 ;
        RECT 539.740 498.710 540.110 498.850 ;
        RECT 539.740 491.630 539.880 498.710 ;
        RECT 539.680 491.310 539.940 491.630 ;
        RECT 541.060 491.310 541.320 491.630 ;
        RECT 541.120 163.870 541.260 491.310 ;
        RECT 541.060 163.550 541.320 163.870 ;
        RECT 1331.800 163.550 1332.060 163.870 ;
        RECT 1331.860 82.870 1332.000 163.550 ;
        RECT 1331.860 82.730 1332.920 82.870 ;
        RECT 1332.780 2.400 1332.920 82.730 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.430 473.520 490.750 473.580 ;
        RECT 494.570 473.520 494.890 473.580 ;
        RECT 490.430 473.380 494.890 473.520 ;
        RECT 490.430 473.320 490.750 473.380 ;
        RECT 494.570 473.320 494.890 473.380 ;
        RECT 493.650 172.280 493.970 172.340 ;
        RECT 690.070 172.280 690.390 172.340 ;
        RECT 493.650 172.140 690.390 172.280 ;
        RECT 493.650 172.080 493.970 172.140 ;
        RECT 690.070 172.080 690.390 172.140 ;
      LAYER via ;
        RECT 490.460 473.320 490.720 473.580 ;
        RECT 494.600 473.320 494.860 473.580 ;
        RECT 493.680 172.080 493.940 172.340 ;
        RECT 690.100 172.080 690.360 172.340 ;
      LAYER met2 ;
        RECT 490.250 500.000 490.530 504.000 ;
        RECT 490.290 499.815 490.430 500.000 ;
        RECT 490.220 499.445 490.500 499.815 ;
        RECT 490.450 497.915 490.730 498.285 ;
        RECT 490.520 473.610 490.660 497.915 ;
        RECT 490.460 473.290 490.720 473.610 ;
        RECT 494.600 473.290 494.860 473.610 ;
        RECT 494.660 448.570 494.800 473.290 ;
        RECT 494.200 448.430 494.800 448.570 ;
        RECT 494.200 420.970 494.340 448.430 ;
        RECT 493.740 420.830 494.340 420.970 ;
        RECT 493.740 172.370 493.880 420.830 ;
        RECT 493.680 172.050 493.940 172.370 ;
        RECT 690.100 172.050 690.360 172.370 ;
        RECT 690.160 82.870 690.300 172.050 ;
        RECT 690.160 82.730 694.440 82.870 ;
        RECT 694.300 2.400 694.440 82.730 ;
        RECT 694.090 -4.800 694.650 2.400 ;
      LAYER via2 ;
        RECT 490.220 499.490 490.500 499.770 ;
        RECT 490.450 497.960 490.730 498.240 ;
      LAYER met3 ;
        RECT 490.195 499.780 490.525 499.795 ;
        RECT 489.520 499.480 490.525 499.780 ;
        RECT 489.520 498.250 489.820 499.480 ;
        RECT 490.195 499.465 490.525 499.480 ;
        RECT 490.425 498.250 490.755 498.265 ;
        RECT 489.520 497.950 490.755 498.250 ;
        RECT 490.425 497.935 490.755 497.950 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 541.950 183.840 542.270 183.900 ;
        RECT 1345.570 183.840 1345.890 183.900 ;
        RECT 541.950 183.700 1345.890 183.840 ;
        RECT 541.950 183.640 542.270 183.700 ;
        RECT 1345.570 183.640 1345.890 183.700 ;
      LAYER via ;
        RECT 541.980 183.640 542.240 183.900 ;
        RECT 1345.600 183.640 1345.860 183.900 ;
      LAYER met2 ;
        RECT 541.310 500.000 541.590 504.000 ;
        RECT 541.350 499.815 541.490 500.000 ;
        RECT 541.280 499.445 541.560 499.815 ;
        RECT 541.510 498.595 541.790 498.965 ;
        RECT 541.580 483.070 541.720 498.595 ;
        RECT 541.580 482.930 542.180 483.070 ;
        RECT 542.040 183.930 542.180 482.930 ;
        RECT 541.980 183.610 542.240 183.930 ;
        RECT 1345.600 183.610 1345.860 183.930 ;
        RECT 1345.660 82.870 1345.800 183.610 ;
        RECT 1345.660 82.730 1350.400 82.870 ;
        RECT 1350.260 2.400 1350.400 82.730 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
      LAYER via2 ;
        RECT 541.280 499.490 541.560 499.770 ;
        RECT 541.510 498.640 541.790 498.920 ;
      LAYER met3 ;
        RECT 541.255 499.465 541.585 499.795 ;
        RECT 541.270 498.945 541.570 499.465 ;
        RECT 541.270 498.630 541.815 498.945 ;
        RECT 541.485 498.615 541.815 498.630 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 542.640 499.160 542.960 499.420 ;
        RECT 542.730 498.340 542.870 499.160 ;
        RECT 542.730 498.200 543.560 498.340 ;
        RECT 541.950 497.660 542.270 497.720 ;
        RECT 543.420 497.660 543.560 498.200 ;
        RECT 541.950 497.520 543.560 497.660 ;
        RECT 541.950 497.460 542.270 497.520 ;
      LAYER via ;
        RECT 542.670 499.160 542.930 499.420 ;
        RECT 541.980 497.460 542.240 497.720 ;
      LAYER met2 ;
        RECT 542.690 500.000 542.970 504.000 ;
        RECT 542.730 499.450 542.870 500.000 ;
        RECT 542.670 499.130 542.930 499.450 ;
        RECT 541.980 497.430 542.240 497.750 ;
        RECT 542.040 491.485 542.180 497.430 ;
        RECT 541.970 491.115 542.250 491.485 ;
        RECT 1366.290 164.035 1366.570 164.405 ;
        RECT 1366.360 1.770 1366.500 164.035 ;
        RECT 1367.990 1.770 1368.550 2.400 ;
        RECT 1366.360 1.630 1368.550 1.770 ;
        RECT 1367.990 -4.800 1368.550 1.630 ;
      LAYER via2 ;
        RECT 541.970 491.160 542.250 491.440 ;
        RECT 1366.290 164.080 1366.570 164.360 ;
      LAYER met3 ;
        RECT 541.230 491.450 541.610 491.460 ;
        RECT 541.945 491.450 542.275 491.465 ;
        RECT 541.230 491.150 542.275 491.450 ;
        RECT 541.230 491.140 541.610 491.150 ;
        RECT 541.945 491.135 542.275 491.150 ;
        RECT 541.230 164.370 541.610 164.380 ;
        RECT 1366.265 164.370 1366.595 164.385 ;
        RECT 541.230 164.070 1366.595 164.370 ;
        RECT 541.230 164.060 541.610 164.070 ;
        RECT 1366.265 164.055 1366.595 164.070 ;
      LAYER via3 ;
        RECT 541.260 491.140 541.580 491.460 ;
        RECT 541.260 164.060 541.580 164.380 ;
      LAYER met4 ;
        RECT 541.255 491.135 541.585 491.465 ;
        RECT 541.270 164.385 541.570 491.135 ;
        RECT 541.255 164.055 541.585 164.385 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 544.020 499.500 544.340 499.760 ;
        RECT 544.110 499.080 544.250 499.500 ;
        RECT 544.110 498.880 544.570 499.080 ;
        RECT 544.250 498.820 544.570 498.880 ;
        RECT 544.250 484.400 544.570 484.460 ;
        RECT 544.250 484.260 591.400 484.400 ;
        RECT 544.250 484.200 544.570 484.260 ;
        RECT 591.260 484.120 591.400 484.260 ;
        RECT 591.170 483.860 591.490 484.120 ;
        RECT 590.710 184.180 591.030 184.240 ;
        RECT 1380.070 184.180 1380.390 184.240 ;
        RECT 590.710 184.040 1380.390 184.180 ;
        RECT 590.710 183.980 591.030 184.040 ;
        RECT 1380.070 183.980 1380.390 184.040 ;
        RECT 1380.070 18.940 1380.390 19.000 ;
        RECT 1383.750 18.940 1384.070 19.000 ;
        RECT 1380.070 18.800 1384.070 18.940 ;
        RECT 1380.070 18.740 1380.390 18.800 ;
        RECT 1383.750 18.740 1384.070 18.800 ;
      LAYER via ;
        RECT 544.050 499.500 544.310 499.760 ;
        RECT 544.280 498.820 544.540 499.080 ;
        RECT 544.280 484.200 544.540 484.460 ;
        RECT 591.200 483.860 591.460 484.120 ;
        RECT 590.740 183.980 591.000 184.240 ;
        RECT 1380.100 183.980 1380.360 184.240 ;
        RECT 1380.100 18.740 1380.360 19.000 ;
        RECT 1383.780 18.740 1384.040 19.000 ;
      LAYER met2 ;
        RECT 544.070 500.000 544.350 504.000 ;
        RECT 544.110 499.790 544.250 500.000 ;
        RECT 544.050 499.470 544.310 499.790 ;
        RECT 544.280 498.790 544.540 499.110 ;
        RECT 544.340 484.490 544.480 498.790 ;
        RECT 544.280 484.170 544.540 484.490 ;
        RECT 591.200 483.830 591.460 484.150 ;
        RECT 591.260 448.570 591.400 483.830 ;
        RECT 590.800 448.430 591.400 448.570 ;
        RECT 590.800 184.270 590.940 448.430 ;
        RECT 590.740 183.950 591.000 184.270 ;
        RECT 1380.100 183.950 1380.360 184.270 ;
        RECT 1380.160 19.030 1380.300 183.950 ;
        RECT 1380.100 18.710 1380.360 19.030 ;
        RECT 1383.780 18.710 1384.040 19.030 ;
        RECT 1383.840 1.770 1383.980 18.710 ;
        RECT 1385.470 1.770 1386.030 2.400 ;
        RECT 1383.840 1.630 1386.030 1.770 ;
        RECT 1385.470 -4.800 1386.030 1.630 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.400 499.160 545.720 499.420 ;
        RECT 545.490 498.000 545.630 499.160 ;
        RECT 546.090 498.000 546.410 498.060 ;
        RECT 545.490 497.860 546.410 498.000 ;
        RECT 546.090 497.800 546.410 497.860 ;
        RECT 545.630 473.520 545.950 473.580 ;
        RECT 547.010 473.520 547.330 473.580 ;
        RECT 545.630 473.380 547.330 473.520 ;
        RECT 545.630 473.320 545.950 473.380 ;
        RECT 547.010 473.320 547.330 473.380 ;
        RECT 547.010 110.400 547.330 110.460 ;
        RECT 1400.770 110.400 1401.090 110.460 ;
        RECT 547.010 110.260 1401.090 110.400 ;
        RECT 547.010 110.200 547.330 110.260 ;
        RECT 1400.770 110.200 1401.090 110.260 ;
      LAYER via ;
        RECT 545.430 499.160 545.690 499.420 ;
        RECT 546.120 497.800 546.380 498.060 ;
        RECT 545.660 473.320 545.920 473.580 ;
        RECT 547.040 473.320 547.300 473.580 ;
        RECT 547.040 110.200 547.300 110.460 ;
        RECT 1400.800 110.200 1401.060 110.460 ;
      LAYER met2 ;
        RECT 545.450 500.000 545.730 504.000 ;
        RECT 545.490 499.450 545.630 500.000 ;
        RECT 545.430 499.130 545.690 499.450 ;
        RECT 546.120 497.770 546.380 498.090 ;
        RECT 546.180 491.540 546.320 497.770 ;
        RECT 545.720 491.400 546.320 491.540 ;
        RECT 545.720 473.610 545.860 491.400 ;
        RECT 545.660 473.290 545.920 473.610 ;
        RECT 547.040 473.290 547.300 473.610 ;
        RECT 547.100 110.490 547.240 473.290 ;
        RECT 547.040 110.170 547.300 110.490 ;
        RECT 1400.800 110.170 1401.060 110.490 ;
        RECT 1400.860 82.870 1401.000 110.170 ;
        RECT 1400.860 82.730 1403.760 82.870 ;
        RECT 1403.620 2.400 1403.760 82.730 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 549.310 183.160 549.630 183.220 ;
        RECT 1421.470 183.160 1421.790 183.220 ;
        RECT 549.310 183.020 1421.790 183.160 ;
        RECT 549.310 182.960 549.630 183.020 ;
        RECT 1421.470 182.960 1421.790 183.020 ;
      LAYER via ;
        RECT 549.340 182.960 549.600 183.220 ;
        RECT 1421.500 182.960 1421.760 183.220 ;
      LAYER met2 ;
        RECT 546.830 500.000 547.110 504.000 ;
        RECT 546.870 499.645 547.010 500.000 ;
        RECT 546.800 499.275 547.080 499.645 ;
        RECT 549.790 497.235 550.070 497.605 ;
        RECT 549.860 420.970 550.000 497.235 ;
        RECT 549.400 420.830 550.000 420.970 ;
        RECT 549.400 183.250 549.540 420.830 ;
        RECT 549.340 182.930 549.600 183.250 ;
        RECT 1421.500 182.930 1421.760 183.250 ;
        RECT 1421.560 2.400 1421.700 182.930 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
      LAYER via2 ;
        RECT 546.800 499.320 547.080 499.600 ;
        RECT 549.790 497.280 550.070 497.560 ;
      LAYER met3 ;
        RECT 546.775 499.295 547.105 499.625 ;
        RECT 546.790 497.570 547.090 499.295 ;
        RECT 549.765 497.570 550.095 497.585 ;
        RECT 546.790 497.270 550.095 497.570 ;
        RECT 549.765 497.255 550.095 497.270 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 548.160 499.500 548.480 499.760 ;
        RECT 548.250 498.400 548.390 499.500 ;
        RECT 547.930 498.200 548.390 498.400 ;
        RECT 547.930 498.140 548.250 498.200 ;
        RECT 547.470 110.060 547.790 110.120 ;
        RECT 1435.270 110.060 1435.590 110.120 ;
        RECT 547.470 109.920 1435.590 110.060 ;
        RECT 547.470 109.860 547.790 109.920 ;
        RECT 1435.270 109.860 1435.590 109.920 ;
      LAYER via ;
        RECT 548.190 499.500 548.450 499.760 ;
        RECT 547.960 498.140 548.220 498.400 ;
        RECT 547.500 109.860 547.760 110.120 ;
        RECT 1435.300 109.860 1435.560 110.120 ;
      LAYER met2 ;
        RECT 548.210 500.000 548.490 504.000 ;
        RECT 548.250 499.790 548.390 500.000 ;
        RECT 548.190 499.470 548.450 499.790 ;
        RECT 547.960 498.110 548.220 498.430 ;
        RECT 548.020 483.070 548.160 498.110 ;
        RECT 547.560 482.930 548.160 483.070 ;
        RECT 547.560 476.170 547.700 482.930 ;
        RECT 547.560 476.030 548.160 476.170 ;
        RECT 548.020 473.010 548.160 476.030 ;
        RECT 547.560 472.870 548.160 473.010 ;
        RECT 547.560 110.150 547.700 472.870 ;
        RECT 547.500 109.830 547.760 110.150 ;
        RECT 1435.300 109.830 1435.560 110.150 ;
        RECT 1435.360 82.870 1435.500 109.830 ;
        RECT 1435.360 82.730 1436.880 82.870 ;
        RECT 1436.740 1.770 1436.880 82.730 ;
        RECT 1438.830 1.770 1439.390 2.400 ;
        RECT 1436.740 1.630 1439.390 1.770 ;
        RECT 1438.830 -4.800 1439.390 1.630 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 549.540 499.500 549.860 499.760 ;
        RECT 549.630 498.000 549.770 499.500 ;
        RECT 551.150 498.000 551.470 498.060 ;
        RECT 549.630 497.860 551.470 498.000 ;
        RECT 551.150 497.800 551.470 497.860 ;
        RECT 591.170 183.500 591.490 183.560 ;
        RECT 1455.970 183.500 1456.290 183.560 ;
        RECT 591.170 183.360 1456.290 183.500 ;
        RECT 591.170 183.300 591.490 183.360 ;
        RECT 1455.970 183.300 1456.290 183.360 ;
      LAYER via ;
        RECT 549.570 499.500 549.830 499.760 ;
        RECT 551.180 497.800 551.440 498.060 ;
        RECT 591.200 183.300 591.460 183.560 ;
        RECT 1456.000 183.300 1456.260 183.560 ;
      LAYER met2 ;
        RECT 549.590 500.000 549.870 504.000 ;
        RECT 549.630 499.790 549.770 500.000 ;
        RECT 549.570 499.470 549.830 499.790 ;
        RECT 551.180 497.770 551.440 498.090 ;
        RECT 551.240 488.765 551.380 497.770 ;
        RECT 551.170 488.395 551.450 488.765 ;
        RECT 593.030 488.395 593.310 488.765 ;
        RECT 593.100 420.970 593.240 488.395 ;
        RECT 591.260 420.830 593.240 420.970 ;
        RECT 591.260 183.590 591.400 420.830 ;
        RECT 591.200 183.270 591.460 183.590 ;
        RECT 1456.000 183.270 1456.260 183.590 ;
        RECT 1456.060 82.870 1456.200 183.270 ;
        RECT 1456.060 82.730 1457.120 82.870 ;
        RECT 1456.980 2.400 1457.120 82.730 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
      LAYER via2 ;
        RECT 551.170 488.440 551.450 488.720 ;
        RECT 593.030 488.440 593.310 488.720 ;
      LAYER met3 ;
        RECT 551.145 488.730 551.475 488.745 ;
        RECT 593.005 488.730 593.335 488.745 ;
        RECT 551.145 488.430 593.335 488.730 ;
        RECT 551.145 488.415 551.475 488.430 ;
        RECT 593.005 488.415 593.335 488.430 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 550.920 499.500 551.240 499.760 ;
        RECT 551.010 499.080 551.150 499.500 ;
        RECT 550.690 498.880 551.150 499.080 ;
        RECT 550.690 498.820 551.010 498.880 ;
      LAYER via ;
        RECT 550.950 499.500 551.210 499.760 ;
        RECT 550.720 498.820 550.980 499.080 ;
      LAYER met2 ;
        RECT 550.970 500.000 551.250 504.000 ;
        RECT 551.010 499.790 551.150 500.000 ;
        RECT 550.950 499.470 551.210 499.790 ;
        RECT 550.720 498.790 550.980 499.110 ;
        RECT 550.780 491.485 550.920 498.790 ;
        RECT 550.710 491.115 550.990 491.485 ;
        RECT 1469.790 100.795 1470.070 101.165 ;
        RECT 1469.860 82.870 1470.000 100.795 ;
        RECT 1469.860 82.730 1474.600 82.870 ;
        RECT 1474.460 2.400 1474.600 82.730 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
      LAYER via2 ;
        RECT 550.710 491.160 550.990 491.440 ;
        RECT 1469.790 100.840 1470.070 101.120 ;
      LAYER met3 ;
        RECT 546.750 491.450 547.130 491.460 ;
        RECT 550.685 491.450 551.015 491.465 ;
        RECT 546.750 491.150 551.015 491.450 ;
        RECT 546.750 491.140 547.130 491.150 ;
        RECT 550.685 491.135 551.015 491.150 ;
        RECT 546.750 101.130 547.130 101.140 ;
        RECT 1469.765 101.130 1470.095 101.145 ;
        RECT 546.750 100.830 1470.095 101.130 ;
        RECT 546.750 100.820 547.130 100.830 ;
        RECT 1469.765 100.815 1470.095 100.830 ;
      LAYER via3 ;
        RECT 546.780 491.140 547.100 491.460 ;
        RECT 546.780 100.820 547.100 101.140 ;
      LAYER met4 ;
        RECT 546.775 491.135 547.105 491.465 ;
        RECT 546.790 101.145 547.090 491.135 ;
        RECT 546.775 100.815 547.105 101.145 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 551.610 471.480 551.930 471.540 ;
        RECT 554.370 471.480 554.690 471.540 ;
        RECT 551.610 471.340 554.690 471.480 ;
        RECT 551.610 471.280 551.930 471.340 ;
        RECT 554.370 471.280 554.690 471.340 ;
        RECT 554.370 102.240 554.690 102.300 ;
        RECT 1490.470 102.240 1490.790 102.300 ;
        RECT 554.370 102.100 1490.790 102.240 ;
        RECT 554.370 102.040 554.690 102.100 ;
        RECT 1490.470 102.040 1490.790 102.100 ;
      LAYER via ;
        RECT 551.640 471.280 551.900 471.540 ;
        RECT 554.400 471.280 554.660 471.540 ;
        RECT 554.400 102.040 554.660 102.300 ;
        RECT 1490.500 102.040 1490.760 102.300 ;
      LAYER met2 ;
        RECT 552.350 500.000 552.630 504.000 ;
        RECT 552.390 499.815 552.530 500.000 ;
        RECT 552.320 499.445 552.600 499.815 ;
        RECT 552.090 497.915 552.370 498.285 ;
        RECT 552.160 473.690 552.300 497.915 ;
        RECT 551.700 473.550 552.300 473.690 ;
        RECT 551.700 471.570 551.840 473.550 ;
        RECT 551.640 471.250 551.900 471.570 ;
        RECT 554.400 471.250 554.660 471.570 ;
        RECT 554.460 102.330 554.600 471.250 ;
        RECT 554.400 102.010 554.660 102.330 ;
        RECT 1490.500 102.010 1490.760 102.330 ;
        RECT 1490.560 1.770 1490.700 102.010 ;
        RECT 1492.190 1.770 1492.750 2.400 ;
        RECT 1490.560 1.630 1492.750 1.770 ;
        RECT 1492.190 -4.800 1492.750 1.630 ;
      LAYER via2 ;
        RECT 552.320 499.490 552.600 499.770 ;
        RECT 552.090 497.960 552.370 498.240 ;
      LAYER met3 ;
        RECT 552.295 499.465 552.625 499.795 ;
        RECT 552.310 498.265 552.610 499.465 ;
        RECT 552.065 497.950 552.610 498.265 ;
        RECT 552.065 497.935 552.395 497.950 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 553.680 500.520 554.000 500.780 ;
        RECT 553.770 500.040 553.910 500.520 ;
        RECT 553.770 499.900 555.290 500.040 ;
        RECT 555.150 498.340 555.290 499.900 ;
        RECT 554.460 498.200 555.290 498.340 ;
        RECT 554.460 496.980 554.600 498.200 ;
        RECT 554.830 496.980 555.150 497.040 ;
        RECT 554.460 496.840 555.150 496.980 ;
        RECT 554.830 496.780 555.150 496.840 ;
        RECT 554.830 109.720 555.150 109.780 ;
        RECT 1504.270 109.720 1504.590 109.780 ;
        RECT 554.830 109.580 1504.590 109.720 ;
        RECT 554.830 109.520 555.150 109.580 ;
        RECT 1504.270 109.520 1504.590 109.580 ;
      LAYER via ;
        RECT 553.710 500.520 553.970 500.780 ;
        RECT 554.860 496.780 555.120 497.040 ;
        RECT 554.860 109.520 555.120 109.780 ;
        RECT 1504.300 109.520 1504.560 109.780 ;
      LAYER met2 ;
        RECT 553.730 500.810 554.010 504.000 ;
        RECT 553.710 500.490 554.010 500.810 ;
        RECT 553.730 500.000 554.010 500.490 ;
        RECT 554.860 496.750 555.120 497.070 ;
        RECT 554.920 109.810 555.060 496.750 ;
        RECT 554.860 109.490 555.120 109.810 ;
        RECT 1504.300 109.490 1504.560 109.810 ;
        RECT 1504.360 82.870 1504.500 109.490 ;
        RECT 1504.360 82.730 1507.720 82.870 ;
        RECT 1507.580 1.770 1507.720 82.730 ;
        RECT 1509.670 1.770 1510.230 2.400 ;
        RECT 1507.580 1.630 1510.230 1.770 ;
        RECT 1509.670 -4.800 1510.230 1.630 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 491.580 501.400 491.900 501.460 ;
        RECT 491.580 501.260 501.700 501.400 ;
        RECT 491.580 501.200 491.900 501.260 ;
        RECT 501.560 498.060 501.700 501.260 ;
        RECT 501.470 497.800 501.790 498.060 ;
        RECT 501.470 486.780 501.790 486.840 ;
        RECT 599.910 486.780 600.230 486.840 ;
        RECT 501.470 486.640 600.230 486.780 ;
        RECT 501.470 486.580 501.790 486.640 ;
        RECT 599.910 486.580 600.230 486.640 ;
        RECT 598.530 181.800 598.850 181.860 ;
        RECT 710.770 181.800 711.090 181.860 ;
        RECT 598.530 181.660 711.090 181.800 ;
        RECT 598.530 181.600 598.850 181.660 ;
        RECT 710.770 181.600 711.090 181.660 ;
      LAYER via ;
        RECT 491.610 501.200 491.870 501.460 ;
        RECT 501.500 497.800 501.760 498.060 ;
        RECT 501.500 486.580 501.760 486.840 ;
        RECT 599.940 486.580 600.200 486.840 ;
        RECT 598.560 181.600 598.820 181.860 ;
        RECT 710.800 181.600 711.060 181.860 ;
      LAYER met2 ;
        RECT 491.630 501.490 491.910 504.000 ;
        RECT 491.610 501.170 491.910 501.490 ;
        RECT 491.630 500.000 491.910 501.170 ;
        RECT 501.500 497.770 501.760 498.090 ;
        RECT 501.560 486.870 501.700 497.770 ;
        RECT 501.500 486.550 501.760 486.870 ;
        RECT 599.940 486.550 600.200 486.870 ;
        RECT 600.000 420.970 600.140 486.550 ;
        RECT 598.620 420.830 600.140 420.970 ;
        RECT 598.620 181.890 598.760 420.830 ;
        RECT 598.560 181.570 598.820 181.890 ;
        RECT 710.800 181.570 711.060 181.890 ;
        RECT 710.860 1.770 711.000 181.570 ;
        RECT 712.030 1.770 712.590 2.400 ;
        RECT 710.860 1.630 712.590 1.770 ;
        RECT 712.030 -4.800 712.590 1.630 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 554.830 497.460 555.150 497.720 ;
        RECT 554.920 497.320 555.060 497.460 ;
        RECT 557.590 497.320 557.910 497.380 ;
        RECT 554.920 497.180 557.910 497.320 ;
        RECT 557.590 497.120 557.910 497.180 ;
        RECT 557.590 483.720 557.910 483.780 ;
        RECT 604.970 483.720 605.290 483.780 ;
        RECT 557.590 483.580 605.290 483.720 ;
        RECT 557.590 483.520 557.910 483.580 ;
        RECT 604.970 483.520 605.290 483.580 ;
        RECT 604.970 193.020 605.290 193.080 ;
        RECT 1524.970 193.020 1525.290 193.080 ;
        RECT 604.970 192.880 1525.290 193.020 ;
        RECT 604.970 192.820 605.290 192.880 ;
        RECT 1524.970 192.820 1525.290 192.880 ;
      LAYER via ;
        RECT 554.860 497.460 555.120 497.720 ;
        RECT 557.620 497.120 557.880 497.380 ;
        RECT 557.620 483.520 557.880 483.780 ;
        RECT 605.000 483.520 605.260 483.780 ;
        RECT 605.000 192.820 605.260 193.080 ;
        RECT 1525.000 192.820 1525.260 193.080 ;
      LAYER met2 ;
        RECT 555.110 500.000 555.390 504.000 ;
        RECT 555.150 498.850 555.290 500.000 ;
        RECT 554.920 498.710 555.290 498.850 ;
        RECT 554.920 497.750 555.060 498.710 ;
        RECT 554.860 497.430 555.120 497.750 ;
        RECT 557.620 497.090 557.880 497.410 ;
        RECT 557.680 483.810 557.820 497.090 ;
        RECT 557.620 483.490 557.880 483.810 ;
        RECT 605.000 483.490 605.260 483.810 ;
        RECT 605.060 193.110 605.200 483.490 ;
        RECT 605.000 192.790 605.260 193.110 ;
        RECT 1525.000 192.790 1525.260 193.110 ;
        RECT 1525.060 82.870 1525.200 192.790 ;
        RECT 1525.060 82.730 1527.960 82.870 ;
        RECT 1527.820 2.400 1527.960 82.730 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1539.230 19.280 1539.550 19.340 ;
        RECT 1545.210 19.280 1545.530 19.340 ;
        RECT 1539.230 19.140 1545.530 19.280 ;
        RECT 1539.230 19.080 1539.550 19.140 ;
        RECT 1545.210 19.080 1545.530 19.140 ;
      LAYER via ;
        RECT 1539.260 19.080 1539.520 19.340 ;
        RECT 1545.240 19.080 1545.500 19.340 ;
      LAYER met2 ;
        RECT 556.490 500.000 556.770 504.000 ;
        RECT 556.530 499.645 556.670 500.000 ;
        RECT 556.460 499.275 556.740 499.645 ;
        RECT 1539.250 106.235 1539.530 106.605 ;
        RECT 1539.320 19.370 1539.460 106.235 ;
        RECT 1539.260 19.050 1539.520 19.370 ;
        RECT 1545.240 19.050 1545.500 19.370 ;
        RECT 1545.300 2.400 1545.440 19.050 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
      LAYER via2 ;
        RECT 556.460 499.320 556.740 499.600 ;
        RECT 1539.250 106.280 1539.530 106.560 ;
      LAYER met3 ;
        RECT 555.030 499.610 555.410 499.620 ;
        RECT 556.435 499.610 556.765 499.625 ;
        RECT 555.030 499.310 556.765 499.610 ;
        RECT 555.030 499.300 555.410 499.310 ;
        RECT 556.435 499.295 556.765 499.310 ;
        RECT 555.030 106.570 555.410 106.580 ;
        RECT 1539.225 106.570 1539.555 106.585 ;
        RECT 555.030 106.270 1539.555 106.570 ;
        RECT 555.030 106.260 555.410 106.270 ;
        RECT 1539.225 106.255 1539.555 106.270 ;
      LAYER via3 ;
        RECT 555.060 499.300 555.380 499.620 ;
        RECT 555.060 106.260 555.380 106.580 ;
      LAYER met4 ;
        RECT 555.055 499.295 555.385 499.625 ;
        RECT 555.070 106.585 555.370 499.295 ;
        RECT 555.055 106.255 555.385 106.585 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 557.820 499.500 558.140 499.760 ;
        RECT 557.910 498.740 558.050 499.500 ;
        RECT 557.910 498.540 558.370 498.740 ;
        RECT 558.050 498.480 558.370 498.540 ;
        RECT 608.190 488.140 608.510 488.200 ;
        RECT 581.140 488.000 608.510 488.140 ;
        RECT 558.050 487.460 558.370 487.520 ;
        RECT 581.140 487.460 581.280 488.000 ;
        RECT 608.190 487.940 608.510 488.000 ;
        RECT 558.050 487.320 581.280 487.460 ;
        RECT 558.050 487.260 558.370 487.320 ;
        RECT 608.190 483.380 608.510 483.440 ;
        RECT 608.190 483.240 611.640 483.380 ;
        RECT 608.190 483.180 608.510 483.240 ;
        RECT 611.500 482.760 611.640 483.240 ;
        RECT 611.410 482.500 611.730 482.760 ;
        RECT 611.870 192.680 612.190 192.740 ;
        RECT 1559.470 192.680 1559.790 192.740 ;
        RECT 611.870 192.540 1559.790 192.680 ;
        RECT 611.870 192.480 612.190 192.540 ;
        RECT 1559.470 192.480 1559.790 192.540 ;
      LAYER via ;
        RECT 557.850 499.500 558.110 499.760 ;
        RECT 558.080 498.480 558.340 498.740 ;
        RECT 558.080 487.260 558.340 487.520 ;
        RECT 608.220 487.940 608.480 488.200 ;
        RECT 608.220 483.180 608.480 483.440 ;
        RECT 611.440 482.500 611.700 482.760 ;
        RECT 611.900 192.480 612.160 192.740 ;
        RECT 1559.500 192.480 1559.760 192.740 ;
      LAYER met2 ;
        RECT 557.870 500.000 558.150 504.000 ;
        RECT 557.910 499.790 558.050 500.000 ;
        RECT 557.850 499.470 558.110 499.790 ;
        RECT 558.080 498.450 558.340 498.770 ;
        RECT 558.140 487.550 558.280 498.450 ;
        RECT 608.220 487.910 608.480 488.230 ;
        RECT 558.080 487.230 558.340 487.550 ;
        RECT 608.280 483.470 608.420 487.910 ;
        RECT 608.220 483.150 608.480 483.470 ;
        RECT 611.440 482.470 611.700 482.790 ;
        RECT 611.500 448.570 611.640 482.470 ;
        RECT 611.500 448.430 612.100 448.570 ;
        RECT 611.960 192.770 612.100 448.430 ;
        RECT 611.900 192.450 612.160 192.770 ;
        RECT 1559.500 192.450 1559.760 192.770 ;
        RECT 1559.560 82.870 1559.700 192.450 ;
        RECT 1559.560 82.730 1561.080 82.870 ;
        RECT 1560.940 1.770 1561.080 82.730 ;
        RECT 1563.030 1.770 1563.590 2.400 ;
        RECT 1560.940 1.630 1563.590 1.770 ;
        RECT 1563.030 -4.800 1563.590 1.630 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.200 499.500 559.520 499.760 ;
        RECT 559.290 499.080 559.430 499.500 ;
        RECT 559.290 498.880 559.750 499.080 ;
        RECT 559.430 498.820 559.750 498.880 ;
        RECT 559.430 472.500 559.750 472.560 ;
        RECT 560.350 472.500 560.670 472.560 ;
        RECT 559.430 472.360 560.670 472.500 ;
        RECT 559.430 472.300 559.750 472.360 ;
        RECT 560.350 472.300 560.670 472.360 ;
        RECT 560.350 109.380 560.670 109.440 ;
        RECT 1580.630 109.380 1580.950 109.440 ;
        RECT 560.350 109.240 1580.950 109.380 ;
        RECT 560.350 109.180 560.670 109.240 ;
        RECT 1580.630 109.180 1580.950 109.240 ;
      LAYER via ;
        RECT 559.230 499.500 559.490 499.760 ;
        RECT 559.460 498.820 559.720 499.080 ;
        RECT 559.460 472.300 559.720 472.560 ;
        RECT 560.380 472.300 560.640 472.560 ;
        RECT 560.380 109.180 560.640 109.440 ;
        RECT 1580.660 109.180 1580.920 109.440 ;
      LAYER met2 ;
        RECT 559.250 500.000 559.530 504.000 ;
        RECT 559.290 499.790 559.430 500.000 ;
        RECT 559.230 499.470 559.490 499.790 ;
        RECT 559.460 498.790 559.720 499.110 ;
        RECT 559.520 472.590 559.660 498.790 ;
        RECT 559.460 472.270 559.720 472.590 ;
        RECT 560.380 472.270 560.640 472.590 ;
        RECT 560.440 109.470 560.580 472.270 ;
        RECT 560.380 109.150 560.640 109.470 ;
        RECT 1580.660 109.150 1580.920 109.470 ;
        RECT 1580.720 82.870 1580.860 109.150 ;
        RECT 1580.720 82.730 1581.320 82.870 ;
        RECT 1581.180 2.400 1581.320 82.730 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 560.810 474.540 561.130 474.600 ;
        RECT 563.110 474.540 563.430 474.600 ;
        RECT 560.810 474.400 563.430 474.540 ;
        RECT 560.810 474.340 561.130 474.400 ;
        RECT 563.110 474.340 563.430 474.400 ;
        RECT 562.650 192.000 562.970 192.060 ;
        RECT 1593.970 192.000 1594.290 192.060 ;
        RECT 562.650 191.860 1594.290 192.000 ;
        RECT 562.650 191.800 562.970 191.860 ;
        RECT 1593.970 191.800 1594.290 191.860 ;
      LAYER via ;
        RECT 560.840 474.340 561.100 474.600 ;
        RECT 563.140 474.340 563.400 474.600 ;
        RECT 562.680 191.800 562.940 192.060 ;
        RECT 1594.000 191.800 1594.260 192.060 ;
      LAYER met2 ;
        RECT 560.630 500.000 560.910 504.000 ;
        RECT 560.670 499.645 560.810 500.000 ;
        RECT 560.600 499.275 560.880 499.645 ;
        RECT 560.830 497.915 561.110 498.285 ;
        RECT 560.900 474.630 561.040 497.915 ;
        RECT 560.840 474.310 561.100 474.630 ;
        RECT 563.140 474.310 563.400 474.630 ;
        RECT 563.200 420.970 563.340 474.310 ;
        RECT 562.740 420.830 563.340 420.970 ;
        RECT 562.740 192.090 562.880 420.830 ;
        RECT 562.680 191.770 562.940 192.090 ;
        RECT 1594.000 191.770 1594.260 192.090 ;
        RECT 1594.060 82.870 1594.200 191.770 ;
        RECT 1594.060 82.730 1598.800 82.870 ;
        RECT 1598.660 2.400 1598.800 82.730 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
      LAYER via2 ;
        RECT 560.600 499.320 560.880 499.600 ;
        RECT 560.830 497.960 561.110 498.240 ;
      LAYER met3 ;
        RECT 560.575 499.295 560.905 499.625 ;
        RECT 560.590 498.265 560.890 499.295 ;
        RECT 560.590 497.950 561.135 498.265 ;
        RECT 560.805 497.935 561.135 497.950 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 562.050 499.900 563.340 500.040 ;
        RECT 562.050 499.760 562.190 499.900 ;
        RECT 561.960 499.500 562.280 499.760 ;
        RECT 562.190 498.680 562.510 498.740 ;
        RECT 563.200 498.680 563.340 499.900 ;
        RECT 562.190 498.540 563.340 498.680 ;
        RECT 562.190 498.480 562.510 498.540 ;
        RECT 562.190 471.280 562.510 471.540 ;
        RECT 562.280 470.520 562.420 471.280 ;
        RECT 562.190 470.260 562.510 470.520 ;
        RECT 562.190 157.660 562.510 157.720 ;
        RECT 1614.670 157.660 1614.990 157.720 ;
        RECT 562.190 157.520 1614.990 157.660 ;
        RECT 562.190 157.460 562.510 157.520 ;
        RECT 1614.670 157.460 1614.990 157.520 ;
      LAYER via ;
        RECT 561.990 499.500 562.250 499.760 ;
        RECT 562.220 498.480 562.480 498.740 ;
        RECT 562.220 471.280 562.480 471.540 ;
        RECT 562.220 470.260 562.480 470.520 ;
        RECT 562.220 157.460 562.480 157.720 ;
        RECT 1614.700 157.460 1614.960 157.720 ;
      LAYER met2 ;
        RECT 562.010 500.000 562.290 504.000 ;
        RECT 562.050 499.790 562.190 500.000 ;
        RECT 561.990 499.470 562.250 499.790 ;
        RECT 562.220 498.450 562.480 498.770 ;
        RECT 562.280 471.570 562.420 498.450 ;
        RECT 562.220 471.250 562.480 471.570 ;
        RECT 562.220 470.230 562.480 470.550 ;
        RECT 562.280 157.750 562.420 470.230 ;
        RECT 562.220 157.430 562.480 157.750 ;
        RECT 1614.700 157.430 1614.960 157.750 ;
        RECT 1614.760 1.770 1614.900 157.430 ;
        RECT 1616.390 1.770 1616.950 2.400 ;
        RECT 1614.760 1.630 1616.950 1.770 ;
        RECT 1616.390 -4.800 1616.950 1.630 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 563.570 487.120 563.890 487.180 ;
        RECT 610.030 487.120 610.350 487.180 ;
        RECT 563.570 486.980 610.350 487.120 ;
        RECT 563.570 486.920 563.890 486.980 ;
        RECT 610.030 486.920 610.350 486.980 ;
        RECT 610.030 482.020 610.350 482.080 ;
        RECT 612.790 482.020 613.110 482.080 ;
        RECT 610.030 481.880 613.110 482.020 ;
        RECT 610.030 481.820 610.350 481.880 ;
        RECT 612.790 481.820 613.110 481.880 ;
        RECT 612.790 192.340 613.110 192.400 ;
        RECT 1628.470 192.340 1628.790 192.400 ;
        RECT 612.790 192.200 1628.790 192.340 ;
        RECT 612.790 192.140 613.110 192.200 ;
        RECT 1628.470 192.140 1628.790 192.200 ;
      LAYER via ;
        RECT 563.600 486.920 563.860 487.180 ;
        RECT 610.060 486.920 610.320 487.180 ;
        RECT 610.060 481.820 610.320 482.080 ;
        RECT 612.820 481.820 613.080 482.080 ;
        RECT 612.820 192.140 613.080 192.400 ;
        RECT 1628.500 192.140 1628.760 192.400 ;
      LAYER met2 ;
        RECT 563.390 500.000 563.670 504.000 ;
        RECT 563.430 498.850 563.570 500.000 ;
        RECT 563.430 498.710 563.800 498.850 ;
        RECT 563.660 487.210 563.800 498.710 ;
        RECT 563.600 486.890 563.860 487.210 ;
        RECT 610.060 486.890 610.320 487.210 ;
        RECT 610.120 482.110 610.260 486.890 ;
        RECT 610.060 481.790 610.320 482.110 ;
        RECT 612.820 481.790 613.080 482.110 ;
        RECT 612.880 192.430 613.020 481.790 ;
        RECT 612.820 192.110 613.080 192.430 ;
        RECT 1628.500 192.110 1628.760 192.430 ;
        RECT 1628.560 82.870 1628.700 192.110 ;
        RECT 1628.560 82.730 1631.920 82.870 ;
        RECT 1631.780 1.770 1631.920 82.730 ;
        RECT 1633.870 1.770 1634.430 2.400 ;
        RECT 1631.780 1.630 1634.430 1.770 ;
        RECT 1633.870 -4.800 1634.430 1.630 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 564.720 499.500 565.040 499.760 ;
        RECT 564.810 499.080 564.950 499.500 ;
        RECT 564.810 498.880 565.270 499.080 ;
        RECT 564.950 498.820 565.270 498.880 ;
      LAYER via ;
        RECT 564.750 499.500 565.010 499.760 ;
        RECT 564.980 498.820 565.240 499.080 ;
      LAYER met2 ;
        RECT 564.770 500.000 565.050 504.000 ;
        RECT 564.810 499.790 564.950 500.000 ;
        RECT 564.750 499.470 565.010 499.790 ;
        RECT 564.980 498.790 565.240 499.110 ;
        RECT 565.040 487.405 565.180 498.790 ;
        RECT 564.970 487.035 565.250 487.405 ;
        RECT 1649.190 163.355 1649.470 163.725 ;
        RECT 1649.260 82.870 1649.400 163.355 ;
        RECT 1649.260 82.730 1652.160 82.870 ;
        RECT 1652.020 2.400 1652.160 82.730 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
      LAYER via2 ;
        RECT 564.970 487.080 565.250 487.360 ;
        RECT 1649.190 163.400 1649.470 163.680 ;
      LAYER met3 ;
        RECT 562.390 487.370 562.770 487.380 ;
        RECT 564.945 487.370 565.275 487.385 ;
        RECT 562.390 487.070 565.275 487.370 ;
        RECT 562.390 487.060 562.770 487.070 ;
        RECT 564.945 487.055 565.275 487.070 ;
        RECT 562.390 163.690 562.770 163.700 ;
        RECT 1649.165 163.690 1649.495 163.705 ;
        RECT 562.390 163.390 1649.495 163.690 ;
        RECT 562.390 163.380 562.770 163.390 ;
        RECT 1649.165 163.375 1649.495 163.390 ;
      LAYER via3 ;
        RECT 562.420 487.060 562.740 487.380 ;
        RECT 562.420 163.380 562.740 163.700 ;
      LAYER met4 ;
        RECT 562.415 487.055 562.745 487.385 ;
        RECT 562.430 163.705 562.730 487.055 ;
        RECT 562.415 163.375 562.745 163.705 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.790 473.520 567.110 473.580 ;
        RECT 570.010 473.520 570.330 473.580 ;
        RECT 566.790 473.380 570.330 473.520 ;
        RECT 566.790 473.320 567.110 473.380 ;
        RECT 570.010 473.320 570.330 473.380 ;
        RECT 569.550 191.660 569.870 191.720 ;
        RECT 1662.970 191.660 1663.290 191.720 ;
        RECT 569.550 191.520 1663.290 191.660 ;
        RECT 569.550 191.460 569.870 191.520 ;
        RECT 1662.970 191.460 1663.290 191.520 ;
        RECT 1662.970 16.900 1663.290 16.960 ;
        RECT 1669.410 16.900 1669.730 16.960 ;
        RECT 1662.970 16.760 1669.730 16.900 ;
        RECT 1662.970 16.700 1663.290 16.760 ;
        RECT 1669.410 16.700 1669.730 16.760 ;
      LAYER via ;
        RECT 566.820 473.320 567.080 473.580 ;
        RECT 570.040 473.320 570.300 473.580 ;
        RECT 569.580 191.460 569.840 191.720 ;
        RECT 1663.000 191.460 1663.260 191.720 ;
        RECT 1663.000 16.700 1663.260 16.960 ;
        RECT 1669.440 16.700 1669.700 16.960 ;
      LAYER met2 ;
        RECT 566.150 500.000 566.430 504.000 ;
        RECT 566.190 499.815 566.330 500.000 ;
        RECT 566.120 499.445 566.400 499.815 ;
        RECT 566.810 491.115 567.090 491.485 ;
        RECT 566.880 473.610 567.020 491.115 ;
        RECT 566.820 473.290 567.080 473.610 ;
        RECT 570.040 473.290 570.300 473.610 ;
        RECT 570.100 448.570 570.240 473.290 ;
        RECT 569.640 448.430 570.240 448.570 ;
        RECT 569.640 191.750 569.780 448.430 ;
        RECT 569.580 191.430 569.840 191.750 ;
        RECT 1663.000 191.430 1663.260 191.750 ;
        RECT 1663.060 16.990 1663.200 191.430 ;
        RECT 1663.000 16.670 1663.260 16.990 ;
        RECT 1669.440 16.670 1669.700 16.990 ;
        RECT 1669.500 2.400 1669.640 16.670 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
      LAYER via2 ;
        RECT 566.120 499.490 566.400 499.770 ;
        RECT 566.810 491.160 567.090 491.440 ;
      LAYER met3 ;
        RECT 566.095 499.620 566.425 499.795 ;
        RECT 566.070 499.610 566.450 499.620 ;
        RECT 566.070 499.310 566.710 499.610 ;
        RECT 566.070 499.300 566.450 499.310 ;
        RECT 566.070 491.450 566.450 491.460 ;
        RECT 566.785 491.450 567.115 491.465 ;
        RECT 566.070 491.150 567.115 491.450 ;
        RECT 566.070 491.140 566.450 491.150 ;
        RECT 566.785 491.135 567.115 491.150 ;
      LAYER via3 ;
        RECT 566.100 499.300 566.420 499.620 ;
        RECT 566.100 491.140 566.420 491.460 ;
      LAYER met4 ;
        RECT 566.095 499.295 566.425 499.625 ;
        RECT 566.110 491.465 566.410 499.295 ;
        RECT 566.095 491.135 566.425 491.465 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 567.480 499.500 567.800 499.760 ;
        RECT 567.570 499.360 567.710 499.500 ;
        RECT 565.500 499.220 567.710 499.360 ;
        RECT 565.500 497.320 565.640 499.220 ;
        RECT 568.630 497.320 568.950 497.380 ;
        RECT 565.500 497.180 568.950 497.320 ;
        RECT 568.630 497.120 568.950 497.180 ;
        RECT 568.630 163.440 568.950 163.500 ;
        RECT 1683.670 163.440 1683.990 163.500 ;
        RECT 568.630 163.300 1683.990 163.440 ;
        RECT 568.630 163.240 568.950 163.300 ;
        RECT 1683.670 163.240 1683.990 163.300 ;
      LAYER via ;
        RECT 567.510 499.500 567.770 499.760 ;
        RECT 568.660 497.120 568.920 497.380 ;
        RECT 568.660 163.240 568.920 163.500 ;
        RECT 1683.700 163.240 1683.960 163.500 ;
      LAYER met2 ;
        RECT 567.530 500.000 567.810 504.000 ;
        RECT 567.570 499.790 567.710 500.000 ;
        RECT 567.510 499.470 567.770 499.790 ;
        RECT 568.660 497.090 568.920 497.410 ;
        RECT 568.720 163.530 568.860 497.090 ;
        RECT 568.660 163.210 568.920 163.530 ;
        RECT 1683.700 163.210 1683.960 163.530 ;
        RECT 1683.760 82.870 1683.900 163.210 ;
        RECT 1683.760 82.730 1685.280 82.870 ;
        RECT 1685.140 1.770 1685.280 82.730 ;
        RECT 1687.230 1.770 1687.790 2.400 ;
        RECT 1685.140 1.630 1687.790 1.770 ;
        RECT 1687.230 -4.800 1687.790 1.630 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 492.960 499.500 493.280 499.760 ;
        RECT 493.050 499.360 493.190 499.500 ;
        RECT 493.050 499.220 493.420 499.360 ;
        RECT 493.280 499.080 493.420 499.220 ;
        RECT 493.190 498.820 493.510 499.080 ;
        RECT 493.190 165.140 493.510 165.200 ;
        RECT 724.570 165.140 724.890 165.200 ;
        RECT 493.190 165.000 724.890 165.140 ;
        RECT 493.190 164.940 493.510 165.000 ;
        RECT 724.570 164.940 724.890 165.000 ;
      LAYER via ;
        RECT 492.990 499.500 493.250 499.760 ;
        RECT 493.220 498.820 493.480 499.080 ;
        RECT 493.220 164.940 493.480 165.200 ;
        RECT 724.600 164.940 724.860 165.200 ;
      LAYER met2 ;
        RECT 493.010 500.000 493.290 504.000 ;
        RECT 493.050 499.790 493.190 500.000 ;
        RECT 492.990 499.470 493.250 499.790 ;
        RECT 493.220 498.790 493.480 499.110 ;
        RECT 493.280 165.230 493.420 498.790 ;
        RECT 493.220 164.910 493.480 165.230 ;
        RECT 724.600 164.910 724.860 165.230 ;
        RECT 724.660 82.870 724.800 164.910 ;
        RECT 724.660 82.730 727.560 82.870 ;
        RECT 727.420 1.770 727.560 82.730 ;
        RECT 729.510 1.770 730.070 2.400 ;
        RECT 727.420 1.630 730.070 1.770 ;
        RECT 729.510 -4.800 730.070 1.630 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 568.860 499.500 569.180 499.760 ;
        RECT 568.950 498.740 569.090 499.500 ;
        RECT 568.950 498.540 569.410 498.740 ;
        RECT 569.090 498.480 569.410 498.540 ;
        RECT 569.090 190.980 569.410 191.040 ;
        RECT 1704.370 190.980 1704.690 191.040 ;
        RECT 569.090 190.840 1704.690 190.980 ;
        RECT 569.090 190.780 569.410 190.840 ;
        RECT 1704.370 190.780 1704.690 190.840 ;
      LAYER via ;
        RECT 568.890 499.500 569.150 499.760 ;
        RECT 569.120 498.480 569.380 498.740 ;
        RECT 569.120 190.780 569.380 191.040 ;
        RECT 1704.400 190.780 1704.660 191.040 ;
      LAYER met2 ;
        RECT 568.910 500.000 569.190 504.000 ;
        RECT 568.950 499.790 569.090 500.000 ;
        RECT 568.890 499.470 569.150 499.790 ;
        RECT 569.120 498.450 569.380 498.770 ;
        RECT 569.180 191.070 569.320 498.450 ;
        RECT 569.120 190.750 569.380 191.070 ;
        RECT 1704.400 190.750 1704.660 191.070 ;
        RECT 1704.460 16.050 1704.600 190.750 ;
        RECT 1704.460 15.910 1705.060 16.050 ;
        RECT 1704.920 2.400 1705.060 15.910 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 570.240 499.500 570.560 499.760 ;
        RECT 570.330 499.080 570.470 499.500 ;
        RECT 570.010 498.880 570.470 499.080 ;
        RECT 570.010 498.820 570.330 498.880 ;
      LAYER via ;
        RECT 570.270 499.500 570.530 499.760 ;
        RECT 570.040 498.820 570.300 499.080 ;
      LAYER met2 ;
        RECT 570.290 500.000 570.570 504.000 ;
        RECT 570.330 499.790 570.470 500.000 ;
        RECT 570.270 499.470 570.530 499.790 ;
        RECT 570.040 498.790 570.300 499.110 ;
        RECT 570.100 491.485 570.240 498.790 ;
        RECT 570.030 491.115 570.310 491.485 ;
        RECT 1718.190 170.155 1718.470 170.525 ;
        RECT 1718.260 82.870 1718.400 170.155 ;
        RECT 1718.260 82.730 1723.000 82.870 ;
        RECT 1722.860 2.400 1723.000 82.730 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
      LAYER via2 ;
        RECT 570.030 491.160 570.310 491.440 ;
        RECT 1718.190 170.200 1718.470 170.480 ;
      LAYER met3 ;
        RECT 567.910 491.450 568.290 491.460 ;
        RECT 570.005 491.450 570.335 491.465 ;
        RECT 567.910 491.150 570.335 491.450 ;
        RECT 567.910 491.140 568.290 491.150 ;
        RECT 570.005 491.135 570.335 491.150 ;
        RECT 567.910 170.490 568.290 170.500 ;
        RECT 1718.165 170.490 1718.495 170.505 ;
        RECT 567.910 170.190 1718.495 170.490 ;
        RECT 567.910 170.180 568.290 170.190 ;
        RECT 1718.165 170.175 1718.495 170.190 ;
      LAYER via3 ;
        RECT 567.940 491.140 568.260 491.460 ;
        RECT 567.940 170.180 568.260 170.500 ;
      LAYER met4 ;
        RECT 567.935 491.135 568.265 491.465 ;
        RECT 567.950 170.505 568.250 491.135 ;
        RECT 567.935 170.175 568.265 170.505 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 571.850 484.740 572.170 484.800 ;
        RECT 618.770 484.740 619.090 484.800 ;
        RECT 571.850 484.600 619.090 484.740 ;
        RECT 571.850 484.540 572.170 484.600 ;
        RECT 618.770 484.540 619.090 484.600 ;
        RECT 619.230 191.320 619.550 191.380 ;
        RECT 1738.870 191.320 1739.190 191.380 ;
        RECT 619.230 191.180 1739.190 191.320 ;
        RECT 619.230 191.120 619.550 191.180 ;
        RECT 1738.870 191.120 1739.190 191.180 ;
      LAYER via ;
        RECT 571.880 484.540 572.140 484.800 ;
        RECT 618.800 484.540 619.060 484.800 ;
        RECT 619.260 191.120 619.520 191.380 ;
        RECT 1738.900 191.120 1739.160 191.380 ;
      LAYER met2 ;
        RECT 571.670 500.000 571.950 504.000 ;
        RECT 571.710 498.680 571.850 500.000 ;
        RECT 571.710 498.540 572.080 498.680 ;
        RECT 571.940 484.830 572.080 498.540 ;
        RECT 571.880 484.510 572.140 484.830 ;
        RECT 618.800 484.510 619.060 484.830 ;
        RECT 618.860 448.570 619.000 484.510 ;
        RECT 618.860 448.430 619.460 448.570 ;
        RECT 619.320 191.410 619.460 448.430 ;
        RECT 619.260 191.090 619.520 191.410 ;
        RECT 1738.900 191.090 1739.160 191.410 ;
        RECT 1738.960 82.870 1739.100 191.090 ;
        RECT 1738.960 82.730 1740.480 82.870 ;
        RECT 1740.340 2.400 1740.480 82.730 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 572.770 472.500 573.090 472.560 ;
        RECT 575.070 472.500 575.390 472.560 ;
        RECT 572.770 472.360 575.390 472.500 ;
        RECT 572.770 472.300 573.090 472.360 ;
        RECT 575.070 472.300 575.390 472.360 ;
        RECT 575.070 116.860 575.390 116.920 ;
        RECT 1752.670 116.860 1752.990 116.920 ;
        RECT 575.070 116.720 1752.990 116.860 ;
        RECT 575.070 116.660 575.390 116.720 ;
        RECT 1752.670 116.660 1752.990 116.720 ;
      LAYER via ;
        RECT 572.800 472.300 573.060 472.560 ;
        RECT 575.100 472.300 575.360 472.560 ;
        RECT 575.100 116.660 575.360 116.920 ;
        RECT 1752.700 116.660 1752.960 116.920 ;
      LAYER met2 ;
        RECT 573.050 500.000 573.330 504.000 ;
        RECT 573.090 498.850 573.230 500.000 ;
        RECT 572.860 498.710 573.230 498.850 ;
        RECT 572.860 472.590 573.000 498.710 ;
        RECT 572.800 472.270 573.060 472.590 ;
        RECT 575.100 472.270 575.360 472.590 ;
        RECT 575.160 116.950 575.300 472.270 ;
        RECT 575.100 116.630 575.360 116.950 ;
        RECT 1752.700 116.630 1752.960 116.950 ;
        RECT 1752.760 82.870 1752.900 116.630 ;
        RECT 1752.760 82.730 1756.120 82.870 ;
        RECT 1755.980 1.770 1756.120 82.730 ;
        RECT 1758.070 1.770 1758.630 2.400 ;
        RECT 1755.980 1.630 1758.630 1.770 ;
        RECT 1758.070 -4.800 1758.630 1.630 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 576.910 488.820 577.230 488.880 ;
        RECT 588.870 488.820 589.190 488.880 ;
        RECT 576.910 488.680 589.190 488.820 ;
        RECT 576.910 488.620 577.230 488.680 ;
        RECT 588.870 488.620 589.190 488.680 ;
        RECT 588.870 487.800 589.190 487.860 ;
        RECT 621.990 487.800 622.310 487.860 ;
        RECT 588.870 487.660 622.310 487.800 ;
        RECT 588.870 487.600 589.190 487.660 ;
        RECT 621.990 487.600 622.310 487.660 ;
        RECT 621.990 483.380 622.310 483.440 ;
        RECT 626.130 483.380 626.450 483.440 ;
        RECT 621.990 483.240 626.450 483.380 ;
        RECT 621.990 483.180 622.310 483.240 ;
        RECT 626.130 483.180 626.450 483.240 ;
        RECT 624.750 190.640 625.070 190.700 ;
        RECT 1773.370 190.640 1773.690 190.700 ;
        RECT 624.750 190.500 1773.690 190.640 ;
        RECT 624.750 190.440 625.070 190.500 ;
        RECT 1773.370 190.440 1773.690 190.500 ;
      LAYER via ;
        RECT 576.940 488.620 577.200 488.880 ;
        RECT 588.900 488.620 589.160 488.880 ;
        RECT 588.900 487.600 589.160 487.860 ;
        RECT 622.020 487.600 622.280 487.860 ;
        RECT 622.020 483.180 622.280 483.440 ;
        RECT 626.160 483.180 626.420 483.440 ;
        RECT 624.780 190.440 625.040 190.700 ;
        RECT 1773.400 190.440 1773.660 190.700 ;
      LAYER met2 ;
        RECT 574.430 500.000 574.710 504.000 ;
        RECT 574.470 499.645 574.610 500.000 ;
        RECT 574.400 499.275 574.680 499.645 ;
        RECT 576.930 498.595 577.210 498.965 ;
        RECT 577.000 488.910 577.140 498.595 ;
        RECT 576.940 488.590 577.200 488.910 ;
        RECT 588.900 488.590 589.160 488.910 ;
        RECT 588.960 487.890 589.100 488.590 ;
        RECT 588.900 487.570 589.160 487.890 ;
        RECT 622.020 487.570 622.280 487.890 ;
        RECT 622.080 483.470 622.220 487.570 ;
        RECT 622.020 483.150 622.280 483.470 ;
        RECT 626.160 483.150 626.420 483.470 ;
        RECT 626.220 448.570 626.360 483.150 ;
        RECT 624.840 448.430 626.360 448.570 ;
        RECT 624.840 190.730 624.980 448.430 ;
        RECT 624.780 190.410 625.040 190.730 ;
        RECT 1773.400 190.410 1773.660 190.730 ;
        RECT 1773.460 82.870 1773.600 190.410 ;
        RECT 1773.460 82.730 1776.360 82.870 ;
        RECT 1776.220 2.400 1776.360 82.730 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
      LAYER via2 ;
        RECT 574.400 499.320 574.680 499.600 ;
        RECT 576.930 498.640 577.210 498.920 ;
      LAYER met3 ;
        RECT 574.375 499.295 574.705 499.625 ;
        RECT 574.390 498.930 574.690 499.295 ;
        RECT 576.905 498.930 577.235 498.945 ;
        RECT 574.390 498.630 577.235 498.930 ;
        RECT 576.905 498.615 577.235 498.630 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.610 116.520 574.930 116.580 ;
        RECT 1787.170 116.520 1787.490 116.580 ;
        RECT 574.610 116.380 1787.490 116.520 ;
        RECT 574.610 116.320 574.930 116.380 ;
        RECT 1787.170 116.320 1787.490 116.380 ;
        RECT 1787.170 16.900 1787.490 16.960 ;
        RECT 1793.610 16.900 1793.930 16.960 ;
        RECT 1787.170 16.760 1793.930 16.900 ;
        RECT 1787.170 16.700 1787.490 16.760 ;
        RECT 1793.610 16.700 1793.930 16.760 ;
      LAYER via ;
        RECT 574.640 116.320 574.900 116.580 ;
        RECT 1787.200 116.320 1787.460 116.580 ;
        RECT 1787.200 16.700 1787.460 16.960 ;
        RECT 1793.640 16.700 1793.900 16.960 ;
      LAYER met2 ;
        RECT 575.810 500.000 576.090 504.000 ;
        RECT 575.850 498.850 575.990 500.000 ;
        RECT 575.620 498.710 575.990 498.850 ;
        RECT 575.620 473.690 575.760 498.710 ;
        RECT 574.700 473.550 575.760 473.690 ;
        RECT 574.700 116.610 574.840 473.550 ;
        RECT 574.640 116.290 574.900 116.610 ;
        RECT 1787.200 116.290 1787.460 116.610 ;
        RECT 1787.260 16.990 1787.400 116.290 ;
        RECT 1787.200 16.670 1787.460 16.990 ;
        RECT 1793.640 16.670 1793.900 16.990 ;
        RECT 1793.700 2.400 1793.840 16.670 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 577.140 499.160 577.460 499.420 ;
        RECT 577.230 497.320 577.370 499.160 ;
        RECT 578.750 497.320 579.070 497.380 ;
        RECT 577.230 497.180 579.070 497.320 ;
        RECT 578.750 497.120 579.070 497.180 ;
        RECT 612.330 190.300 612.650 190.360 ;
        RECT 1807.870 190.300 1808.190 190.360 ;
        RECT 612.330 190.160 1808.190 190.300 ;
        RECT 612.330 190.100 612.650 190.160 ;
        RECT 1807.870 190.100 1808.190 190.160 ;
      LAYER via ;
        RECT 577.170 499.160 577.430 499.420 ;
        RECT 578.780 497.120 579.040 497.380 ;
        RECT 612.360 190.100 612.620 190.360 ;
        RECT 1807.900 190.100 1808.160 190.360 ;
      LAYER met2 ;
        RECT 577.190 500.000 577.470 504.000 ;
        RECT 577.230 499.450 577.370 500.000 ;
        RECT 577.170 499.130 577.430 499.450 ;
        RECT 578.780 497.090 579.040 497.410 ;
        RECT 578.840 487.405 578.980 497.090 ;
        RECT 578.770 487.035 579.050 487.405 ;
        RECT 613.730 487.035 614.010 487.405 ;
        RECT 613.800 482.530 613.940 487.035 ;
        RECT 612.420 482.390 613.940 482.530 ;
        RECT 612.420 190.390 612.560 482.390 ;
        RECT 612.360 190.070 612.620 190.390 ;
        RECT 1807.900 190.070 1808.160 190.390 ;
        RECT 1807.960 82.870 1808.100 190.070 ;
        RECT 1807.960 82.730 1809.480 82.870 ;
        RECT 1809.340 1.770 1809.480 82.730 ;
        RECT 1811.430 1.770 1811.990 2.400 ;
        RECT 1809.340 1.630 1811.990 1.770 ;
        RECT 1811.430 -4.800 1811.990 1.630 ;
      LAYER via2 ;
        RECT 578.770 487.080 579.050 487.360 ;
        RECT 613.730 487.080 614.010 487.360 ;
      LAYER met3 ;
        RECT 578.745 487.370 579.075 487.385 ;
        RECT 613.705 487.370 614.035 487.385 ;
        RECT 578.745 487.070 614.035 487.370 ;
        RECT 578.745 487.055 579.075 487.070 ;
        RECT 613.705 487.055 614.035 487.070 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.570 500.000 578.850 504.000 ;
        RECT 578.610 498.000 578.750 500.000 ;
        RECT 578.380 497.860 578.750 498.000 ;
        RECT 578.380 484.005 578.520 497.860 ;
        RECT 578.310 483.635 578.590 484.005 ;
        RECT 1828.590 113.035 1828.870 113.405 ;
        RECT 1828.660 16.050 1828.800 113.035 ;
        RECT 1828.660 15.910 1829.260 16.050 ;
        RECT 1829.120 2.400 1829.260 15.910 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
      LAYER via2 ;
        RECT 578.310 483.680 578.590 483.960 ;
        RECT 1828.590 113.080 1828.870 113.360 ;
      LAYER met3 ;
        RECT 577.110 483.970 577.490 483.980 ;
        RECT 578.285 483.970 578.615 483.985 ;
        RECT 577.110 483.670 578.615 483.970 ;
        RECT 577.110 483.660 577.490 483.670 ;
        RECT 578.285 483.655 578.615 483.670 ;
        RECT 577.110 113.370 577.490 113.380 ;
        RECT 1828.565 113.370 1828.895 113.385 ;
        RECT 577.110 113.070 1828.895 113.370 ;
        RECT 577.110 113.060 577.490 113.070 ;
        RECT 1828.565 113.055 1828.895 113.070 ;
      LAYER via3 ;
        RECT 577.140 483.660 577.460 483.980 ;
        RECT 577.140 113.060 577.460 113.380 ;
      LAYER met4 ;
        RECT 577.135 483.655 577.465 483.985 ;
        RECT 577.150 113.385 577.450 483.655 ;
        RECT 577.135 113.055 577.465 113.385 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.130 495.280 580.450 495.340 ;
        RECT 604.510 495.280 604.830 495.340 ;
        RECT 580.130 495.140 604.830 495.280 ;
        RECT 580.130 495.080 580.450 495.140 ;
        RECT 604.510 495.080 604.830 495.140 ;
        RECT 604.510 486.780 604.830 486.840 ;
        RECT 627.510 486.780 627.830 486.840 ;
        RECT 604.510 486.640 627.830 486.780 ;
        RECT 604.510 486.580 604.830 486.640 ;
        RECT 627.510 486.580 627.830 486.640 ;
        RECT 626.590 189.960 626.910 190.020 ;
        RECT 1842.370 189.960 1842.690 190.020 ;
        RECT 626.590 189.820 1842.690 189.960 ;
        RECT 626.590 189.760 626.910 189.820 ;
        RECT 1842.370 189.760 1842.690 189.820 ;
      LAYER via ;
        RECT 580.160 495.080 580.420 495.340 ;
        RECT 604.540 495.080 604.800 495.340 ;
        RECT 604.540 486.580 604.800 486.840 ;
        RECT 627.540 486.580 627.800 486.840 ;
        RECT 626.620 189.760 626.880 190.020 ;
        RECT 1842.400 189.760 1842.660 190.020 ;
      LAYER met2 ;
        RECT 579.950 500.000 580.230 504.000 ;
        RECT 579.990 499.020 580.130 500.000 ;
        RECT 579.990 498.880 580.360 499.020 ;
        RECT 580.220 495.370 580.360 498.880 ;
        RECT 580.160 495.050 580.420 495.370 ;
        RECT 604.540 495.050 604.800 495.370 ;
        RECT 604.600 486.870 604.740 495.050 ;
        RECT 604.540 486.550 604.800 486.870 ;
        RECT 627.540 486.550 627.800 486.870 ;
        RECT 627.600 448.570 627.740 486.550 ;
        RECT 626.680 448.430 627.740 448.570 ;
        RECT 626.680 190.050 626.820 448.430 ;
        RECT 626.620 189.730 626.880 190.050 ;
        RECT 1842.400 189.730 1842.660 190.050 ;
        RECT 1842.460 82.870 1842.600 189.730 ;
        RECT 1842.460 82.730 1847.200 82.870 ;
        RECT 1847.060 2.400 1847.200 82.730 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 581.280 500.180 581.600 500.440 ;
        RECT 581.370 497.660 581.510 500.180 ;
        RECT 583.350 497.660 583.670 497.720 ;
        RECT 581.370 497.520 583.670 497.660 ;
        RECT 583.350 497.460 583.670 497.520 ;
        RECT 582.890 171.260 583.210 171.320 ;
        RECT 1863.070 171.260 1863.390 171.320 ;
        RECT 582.890 171.120 1863.390 171.260 ;
        RECT 582.890 171.060 583.210 171.120 ;
        RECT 1863.070 171.060 1863.390 171.120 ;
      LAYER via ;
        RECT 581.310 500.180 581.570 500.440 ;
        RECT 583.380 497.460 583.640 497.720 ;
        RECT 582.920 171.060 583.180 171.320 ;
        RECT 1863.100 171.060 1863.360 171.320 ;
      LAYER met2 ;
        RECT 581.330 500.470 581.610 504.000 ;
        RECT 581.310 500.150 581.610 500.470 ;
        RECT 581.330 500.000 581.610 500.150 ;
        RECT 583.380 497.430 583.640 497.750 ;
        RECT 583.440 420.970 583.580 497.430 ;
        RECT 582.980 420.830 583.580 420.970 ;
        RECT 582.980 171.350 583.120 420.830 ;
        RECT 582.920 171.030 583.180 171.350 ;
        RECT 1863.100 171.030 1863.360 171.350 ;
        RECT 1863.160 82.870 1863.300 171.030 ;
        RECT 1863.160 82.730 1864.680 82.870 ;
        RECT 1864.540 2.400 1864.680 82.730 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 491.440 499.900 494.570 500.040 ;
        RECT 491.440 498.740 491.580 499.900 ;
        RECT 494.430 499.760 494.570 499.900 ;
        RECT 494.340 499.500 494.660 499.760 ;
        RECT 491.350 498.480 491.670 498.740 ;
      LAYER via ;
        RECT 494.370 499.500 494.630 499.760 ;
        RECT 491.380 498.480 491.640 498.740 ;
      LAYER met2 ;
        RECT 494.390 500.000 494.670 504.000 ;
        RECT 494.430 499.790 494.570 500.000 ;
        RECT 494.370 499.470 494.630 499.790 ;
        RECT 491.380 498.450 491.640 498.770 ;
        RECT 491.440 487.405 491.580 498.450 ;
        RECT 491.370 487.035 491.650 487.405 ;
        RECT 745.290 114.395 745.570 114.765 ;
        RECT 745.360 82.870 745.500 114.395 ;
        RECT 745.360 82.730 747.800 82.870 ;
        RECT 747.660 2.400 747.800 82.730 ;
        RECT 747.450 -4.800 748.010 2.400 ;
      LAYER via2 ;
        RECT 491.370 487.080 491.650 487.360 ;
        RECT 745.290 114.440 745.570 114.720 ;
      LAYER met3 ;
        RECT 491.345 487.370 491.675 487.385 ;
        RECT 495.230 487.370 495.610 487.380 ;
        RECT 491.345 487.070 495.610 487.370 ;
        RECT 491.345 487.055 491.675 487.070 ;
        RECT 495.230 487.060 495.610 487.070 ;
        RECT 495.230 114.730 495.610 114.740 ;
        RECT 745.265 114.730 745.595 114.745 ;
        RECT 495.230 114.430 745.595 114.730 ;
        RECT 495.230 114.420 495.610 114.430 ;
        RECT 745.265 114.415 745.595 114.430 ;
      LAYER via3 ;
        RECT 495.260 487.060 495.580 487.380 ;
        RECT 495.260 114.420 495.580 114.740 ;
      LAYER met4 ;
        RECT 495.255 487.055 495.585 487.385 ;
        RECT 495.270 114.745 495.570 487.055 ;
        RECT 495.255 114.415 495.585 114.745 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 582.430 498.340 582.750 498.400 ;
        RECT 584.730 498.340 585.050 498.400 ;
        RECT 582.430 498.200 585.050 498.340 ;
        RECT 582.430 498.140 582.750 498.200 ;
        RECT 584.730 498.140 585.050 498.200 ;
        RECT 584.730 490.860 585.050 490.920 ;
        RECT 605.890 490.860 606.210 490.920 ;
        RECT 584.730 490.720 606.210 490.860 ;
        RECT 584.730 490.660 585.050 490.720 ;
        RECT 605.890 490.660 606.210 490.720 ;
        RECT 605.430 382.740 605.750 382.800 ;
        RECT 1876.870 382.740 1877.190 382.800 ;
        RECT 605.430 382.600 1877.190 382.740 ;
        RECT 605.430 382.540 605.750 382.600 ;
        RECT 1876.870 382.540 1877.190 382.600 ;
      LAYER via ;
        RECT 582.460 498.140 582.720 498.400 ;
        RECT 584.760 498.140 585.020 498.400 ;
        RECT 584.760 490.660 585.020 490.920 ;
        RECT 605.920 490.660 606.180 490.920 ;
        RECT 605.460 382.540 605.720 382.800 ;
        RECT 1876.900 382.540 1877.160 382.800 ;
      LAYER met2 ;
        RECT 582.710 500.000 582.990 504.000 ;
        RECT 582.750 499.020 582.890 500.000 ;
        RECT 582.520 498.880 582.890 499.020 ;
        RECT 582.520 498.430 582.660 498.880 ;
        RECT 582.460 498.110 582.720 498.430 ;
        RECT 584.760 498.110 585.020 498.430 ;
        RECT 584.820 490.950 584.960 498.110 ;
        RECT 584.760 490.630 585.020 490.950 ;
        RECT 605.920 490.630 606.180 490.950 ;
        RECT 605.980 448.570 606.120 490.630 ;
        RECT 605.520 448.430 606.120 448.570 ;
        RECT 605.520 382.830 605.660 448.430 ;
        RECT 605.460 382.510 605.720 382.830 ;
        RECT 1876.900 382.510 1877.160 382.830 ;
        RECT 1876.960 82.870 1877.100 382.510 ;
        RECT 1876.960 82.730 1880.320 82.870 ;
        RECT 1880.180 1.770 1880.320 82.730 ;
        RECT 1882.270 1.770 1882.830 2.400 ;
        RECT 1880.180 1.630 1882.830 1.770 ;
        RECT 1882.270 -4.800 1882.830 1.630 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 584.040 499.500 584.360 499.760 ;
        RECT 584.130 499.080 584.270 499.500 ;
        RECT 583.810 498.880 584.270 499.080 ;
        RECT 583.810 498.820 584.130 498.880 ;
        RECT 582.890 490.860 583.210 490.920 ;
        RECT 583.810 490.860 584.130 490.920 ;
        RECT 582.890 490.720 584.130 490.860 ;
        RECT 582.890 490.660 583.210 490.720 ;
        RECT 583.810 490.660 584.130 490.720 ;
        RECT 582.430 170.920 582.750 170.980 ;
        RECT 1897.570 170.920 1897.890 170.980 ;
        RECT 582.430 170.780 1897.890 170.920 ;
        RECT 582.430 170.720 582.750 170.780 ;
        RECT 1897.570 170.720 1897.890 170.780 ;
      LAYER via ;
        RECT 584.070 499.500 584.330 499.760 ;
        RECT 583.840 498.820 584.100 499.080 ;
        RECT 582.920 490.660 583.180 490.920 ;
        RECT 583.840 490.660 584.100 490.920 ;
        RECT 582.460 170.720 582.720 170.980 ;
        RECT 1897.600 170.720 1897.860 170.980 ;
      LAYER met2 ;
        RECT 584.090 500.000 584.370 504.000 ;
        RECT 584.130 499.790 584.270 500.000 ;
        RECT 584.070 499.470 584.330 499.790 ;
        RECT 583.840 498.790 584.100 499.110 ;
        RECT 583.900 490.950 584.040 498.790 ;
        RECT 582.920 490.630 583.180 490.950 ;
        RECT 583.840 490.630 584.100 490.950 ;
        RECT 582.980 448.570 583.120 490.630 ;
        RECT 582.520 448.430 583.120 448.570 ;
        RECT 582.520 171.010 582.660 448.430 ;
        RECT 582.460 170.690 582.720 171.010 ;
        RECT 1897.600 170.690 1897.860 171.010 ;
        RECT 1897.660 1.770 1897.800 170.690 ;
        RECT 1899.750 1.770 1900.310 2.400 ;
        RECT 1897.660 1.630 1900.310 1.770 ;
        RECT 1899.750 -4.800 1900.310 1.630 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1911.370 16.900 1911.690 16.960 ;
        RECT 1917.810 16.900 1918.130 16.960 ;
        RECT 1911.370 16.760 1918.130 16.900 ;
        RECT 1911.370 16.700 1911.690 16.760 ;
        RECT 1917.810 16.700 1918.130 16.760 ;
      LAYER via ;
        RECT 1911.400 16.700 1911.660 16.960 ;
        RECT 1917.840 16.700 1918.100 16.960 ;
      LAYER met2 ;
        RECT 585.470 500.000 585.750 504.000 ;
        RECT 585.510 498.680 585.650 500.000 ;
        RECT 585.280 498.540 585.650 498.680 ;
        RECT 585.280 492.165 585.420 498.540 ;
        RECT 585.210 491.795 585.490 492.165 ;
        RECT 1911.390 162.675 1911.670 163.045 ;
        RECT 1911.460 16.990 1911.600 162.675 ;
        RECT 1911.400 16.670 1911.660 16.990 ;
        RECT 1917.840 16.670 1918.100 16.990 ;
        RECT 1917.900 2.400 1918.040 16.670 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
      LAYER via2 ;
        RECT 585.210 491.840 585.490 492.120 ;
        RECT 1911.390 162.720 1911.670 163.000 ;
      LAYER met3 ;
        RECT 582.630 492.130 583.010 492.140 ;
        RECT 585.185 492.130 585.515 492.145 ;
        RECT 582.630 491.830 585.515 492.130 ;
        RECT 582.630 491.820 583.010 491.830 ;
        RECT 585.185 491.815 585.515 491.830 ;
        RECT 582.630 163.010 583.010 163.020 ;
        RECT 1911.365 163.010 1911.695 163.025 ;
        RECT 582.630 162.710 1911.695 163.010 ;
        RECT 582.630 162.700 583.010 162.710 ;
        RECT 1911.365 162.695 1911.695 162.710 ;
      LAYER via3 ;
        RECT 582.660 491.820 582.980 492.140 ;
        RECT 582.660 162.700 582.980 163.020 ;
      LAYER met4 ;
        RECT 582.655 491.815 582.985 492.145 ;
        RECT 582.670 163.025 582.970 491.815 ;
        RECT 582.655 162.695 582.985 163.025 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.800 499.700 587.120 499.760 ;
        RECT 586.800 499.500 587.260 499.700 ;
        RECT 587.120 497.660 587.260 499.500 ;
        RECT 590.250 497.660 590.570 497.720 ;
        RECT 587.120 497.520 590.570 497.660 ;
        RECT 590.250 497.460 590.570 497.520 ;
        RECT 589.790 170.580 590.110 170.640 ;
        RECT 1932.070 170.580 1932.390 170.640 ;
        RECT 589.790 170.440 1932.390 170.580 ;
        RECT 589.790 170.380 590.110 170.440 ;
        RECT 1932.070 170.380 1932.390 170.440 ;
      LAYER via ;
        RECT 586.830 499.500 587.090 499.760 ;
        RECT 590.280 497.460 590.540 497.720 ;
        RECT 589.820 170.380 590.080 170.640 ;
        RECT 1932.100 170.380 1932.360 170.640 ;
      LAYER met2 ;
        RECT 586.850 500.000 587.130 504.000 ;
        RECT 586.890 499.790 587.030 500.000 ;
        RECT 586.830 499.470 587.090 499.790 ;
        RECT 590.280 497.430 590.540 497.750 ;
        RECT 590.340 492.730 590.480 497.430 ;
        RECT 590.340 492.590 590.940 492.730 ;
        RECT 590.800 473.010 590.940 492.590 ;
        RECT 589.880 472.870 590.940 473.010 ;
        RECT 589.880 170.670 590.020 472.870 ;
        RECT 589.820 170.350 590.080 170.670 ;
        RECT 1932.100 170.350 1932.360 170.670 ;
        RECT 1932.160 82.870 1932.300 170.350 ;
        RECT 1932.160 82.730 1933.680 82.870 ;
        RECT 1933.540 1.770 1933.680 82.730 ;
        RECT 1935.630 1.770 1936.190 2.400 ;
        RECT 1933.540 1.630 1936.190 1.770 ;
        RECT 1935.630 -4.800 1936.190 1.630 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 588.180 499.500 588.500 499.760 ;
        RECT 588.270 499.080 588.410 499.500 ;
        RECT 587.950 498.880 588.410 499.080 ;
        RECT 587.950 498.820 588.270 498.880 ;
        RECT 587.950 494.600 588.270 494.660 ;
        RECT 594.850 494.600 595.170 494.660 ;
        RECT 587.950 494.460 595.170 494.600 ;
        RECT 587.950 494.400 588.270 494.460 ;
        RECT 594.850 494.400 595.170 494.460 ;
        RECT 594.850 485.080 595.170 485.140 ;
        RECT 627.970 485.080 628.290 485.140 ;
        RECT 594.850 484.940 628.290 485.080 ;
        RECT 594.850 484.880 595.170 484.940 ;
        RECT 627.970 484.880 628.290 484.940 ;
        RECT 627.970 483.380 628.290 483.440 ;
        RECT 633.030 483.380 633.350 483.440 ;
        RECT 627.970 483.240 633.350 483.380 ;
        RECT 627.970 483.180 628.290 483.240 ;
        RECT 633.030 483.180 633.350 483.240 ;
        RECT 633.030 108.700 633.350 108.760 ;
        RECT 1953.230 108.700 1953.550 108.760 ;
        RECT 633.030 108.560 1953.550 108.700 ;
        RECT 633.030 108.500 633.350 108.560 ;
        RECT 1953.230 108.500 1953.550 108.560 ;
      LAYER via ;
        RECT 588.210 499.500 588.470 499.760 ;
        RECT 587.980 498.820 588.240 499.080 ;
        RECT 587.980 494.400 588.240 494.660 ;
        RECT 594.880 494.400 595.140 494.660 ;
        RECT 594.880 484.880 595.140 485.140 ;
        RECT 628.000 484.880 628.260 485.140 ;
        RECT 628.000 483.180 628.260 483.440 ;
        RECT 633.060 483.180 633.320 483.440 ;
        RECT 633.060 108.500 633.320 108.760 ;
        RECT 1953.260 108.500 1953.520 108.760 ;
      LAYER met2 ;
        RECT 588.230 500.000 588.510 504.000 ;
        RECT 588.270 499.790 588.410 500.000 ;
        RECT 588.210 499.470 588.470 499.790 ;
        RECT 587.980 498.790 588.240 499.110 ;
        RECT 588.040 494.690 588.180 498.790 ;
        RECT 587.980 494.370 588.240 494.690 ;
        RECT 594.880 494.370 595.140 494.690 ;
        RECT 594.940 485.170 595.080 494.370 ;
        RECT 594.880 484.850 595.140 485.170 ;
        RECT 628.000 484.850 628.260 485.170 ;
        RECT 628.060 483.470 628.200 484.850 ;
        RECT 628.000 483.150 628.260 483.470 ;
        RECT 633.060 483.150 633.320 483.470 ;
        RECT 633.120 108.790 633.260 483.150 ;
        RECT 633.060 108.470 633.320 108.790 ;
        RECT 1953.260 108.470 1953.520 108.790 ;
        RECT 1953.320 2.400 1953.460 108.470 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 589.560 499.500 589.880 499.760 ;
        RECT 589.650 498.740 589.790 499.500 ;
        RECT 589.330 498.540 589.790 498.740 ;
        RECT 589.330 498.480 589.650 498.540 ;
        RECT 589.330 170.240 589.650 170.300 ;
        RECT 1966.570 170.240 1966.890 170.300 ;
        RECT 589.330 170.100 1966.890 170.240 ;
        RECT 589.330 170.040 589.650 170.100 ;
        RECT 1966.570 170.040 1966.890 170.100 ;
      LAYER via ;
        RECT 589.590 499.500 589.850 499.760 ;
        RECT 589.360 498.480 589.620 498.740 ;
        RECT 589.360 170.040 589.620 170.300 ;
        RECT 1966.600 170.040 1966.860 170.300 ;
      LAYER met2 ;
        RECT 589.610 500.000 589.890 504.000 ;
        RECT 589.650 499.790 589.790 500.000 ;
        RECT 589.590 499.470 589.850 499.790 ;
        RECT 589.360 498.450 589.620 498.770 ;
        RECT 589.420 170.330 589.560 498.450 ;
        RECT 589.360 170.010 589.620 170.330 ;
        RECT 1966.600 170.010 1966.860 170.330 ;
        RECT 1966.660 82.870 1966.800 170.010 ;
        RECT 1966.660 82.730 1971.400 82.870 ;
        RECT 1971.260 2.400 1971.400 82.730 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 590.940 499.500 591.260 499.760 ;
        RECT 591.030 498.680 591.170 499.500 ;
        RECT 591.030 498.540 591.860 498.680 ;
        RECT 591.720 498.400 591.860 498.540 ;
        RECT 591.630 498.140 591.950 498.400 ;
        RECT 591.630 494.260 591.950 494.320 ;
        RECT 1987.270 494.260 1987.590 494.320 ;
        RECT 591.630 494.120 1987.590 494.260 ;
        RECT 591.630 494.060 591.950 494.120 ;
        RECT 1987.270 494.060 1987.590 494.120 ;
      LAYER via ;
        RECT 590.970 499.500 591.230 499.760 ;
        RECT 591.660 498.140 591.920 498.400 ;
        RECT 591.660 494.060 591.920 494.320 ;
        RECT 1987.300 494.060 1987.560 494.320 ;
      LAYER met2 ;
        RECT 590.990 500.000 591.270 504.000 ;
        RECT 591.030 499.790 591.170 500.000 ;
        RECT 590.970 499.470 591.230 499.790 ;
        RECT 591.660 498.110 591.920 498.430 ;
        RECT 591.720 494.350 591.860 498.110 ;
        RECT 591.660 494.030 591.920 494.350 ;
        RECT 1987.300 494.030 1987.560 494.350 ;
        RECT 1987.360 82.870 1987.500 494.030 ;
        RECT 1987.360 82.730 1988.880 82.870 ;
        RECT 1988.740 2.400 1988.880 82.730 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 592.320 499.160 592.640 499.420 ;
        RECT 592.410 498.400 592.550 499.160 ;
        RECT 592.090 498.200 592.550 498.400 ;
        RECT 592.090 498.140 592.410 498.200 ;
      LAYER via ;
        RECT 592.350 499.160 592.610 499.420 ;
        RECT 592.120 498.140 592.380 498.400 ;
      LAYER met2 ;
        RECT 592.370 500.000 592.650 504.000 ;
        RECT 592.410 499.450 592.550 500.000 ;
        RECT 592.350 499.130 592.610 499.450 ;
        RECT 592.120 498.110 592.380 498.430 ;
        RECT 592.180 492.845 592.320 498.110 ;
        RECT 592.110 492.475 592.390 492.845 ;
        RECT 2001.090 169.475 2001.370 169.845 ;
        RECT 2001.160 82.870 2001.300 169.475 ;
        RECT 2001.160 82.730 2004.520 82.870 ;
        RECT 2004.380 1.770 2004.520 82.730 ;
        RECT 2006.470 1.770 2007.030 2.400 ;
        RECT 2004.380 1.630 2007.030 1.770 ;
        RECT 2006.470 -4.800 2007.030 1.630 ;
      LAYER via2 ;
        RECT 592.110 492.520 592.390 492.800 ;
        RECT 2001.090 169.520 2001.370 169.800 ;
      LAYER met3 ;
        RECT 589.990 492.810 590.370 492.820 ;
        RECT 592.085 492.810 592.415 492.825 ;
        RECT 589.990 492.510 592.415 492.810 ;
        RECT 589.990 492.500 590.370 492.510 ;
        RECT 592.085 492.495 592.415 492.510 ;
        RECT 589.990 169.810 590.370 169.820 ;
        RECT 2001.065 169.810 2001.395 169.825 ;
        RECT 589.990 169.510 2001.395 169.810 ;
        RECT 589.990 169.500 590.370 169.510 ;
        RECT 2001.065 169.495 2001.395 169.510 ;
      LAYER via3 ;
        RECT 590.020 492.500 590.340 492.820 ;
        RECT 590.020 169.500 590.340 169.820 ;
      LAYER met4 ;
        RECT 590.015 492.495 590.345 492.825 ;
        RECT 590.030 169.825 590.330 492.495 ;
        RECT 590.015 169.495 590.345 169.825 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.700 499.360 594.020 499.420 ;
        RECT 593.700 499.220 595.080 499.360 ;
        RECT 593.700 499.160 594.020 499.220 ;
        RECT 594.940 498.060 595.080 499.220 ;
        RECT 594.850 497.800 595.170 498.060 ;
        RECT 641.310 488.820 641.630 488.880 ;
        RECT 1376.390 488.820 1376.710 488.880 ;
        RECT 641.310 488.680 1376.710 488.820 ;
        RECT 641.310 488.620 641.630 488.680 ;
        RECT 1376.390 488.620 1376.710 488.680 ;
        RECT 602.210 487.460 602.530 487.520 ;
        RECT 641.310 487.460 641.630 487.520 ;
        RECT 602.210 487.320 641.630 487.460 ;
        RECT 602.210 487.260 602.530 487.320 ;
        RECT 641.310 487.260 641.630 487.320 ;
        RECT 1376.390 19.280 1376.710 19.340 ;
        RECT 1376.390 19.140 1386.970 19.280 ;
        RECT 1376.390 19.080 1376.710 19.140 ;
        RECT 1386.830 18.940 1386.970 19.140 ;
        RECT 2024.070 18.940 2024.390 19.000 ;
        RECT 1386.830 18.800 2024.390 18.940 ;
        RECT 2024.070 18.740 2024.390 18.800 ;
      LAYER via ;
        RECT 593.730 499.160 593.990 499.420 ;
        RECT 594.880 497.800 595.140 498.060 ;
        RECT 641.340 488.620 641.600 488.880 ;
        RECT 1376.420 488.620 1376.680 488.880 ;
        RECT 602.240 487.260 602.500 487.520 ;
        RECT 641.340 487.260 641.600 487.520 ;
        RECT 1376.420 19.080 1376.680 19.340 ;
        RECT 2024.100 18.740 2024.360 19.000 ;
      LAYER met2 ;
        RECT 593.750 500.000 594.030 504.000 ;
        RECT 593.790 499.450 593.930 500.000 ;
        RECT 593.730 499.130 593.990 499.450 ;
        RECT 594.880 497.770 595.140 498.090 ;
        RECT 594.940 496.925 595.080 497.770 ;
        RECT 594.870 496.555 595.150 496.925 ;
        RECT 602.230 495.875 602.510 496.245 ;
        RECT 602.300 487.550 602.440 495.875 ;
        RECT 641.340 488.590 641.600 488.910 ;
        RECT 1376.420 488.590 1376.680 488.910 ;
        RECT 641.400 487.550 641.540 488.590 ;
        RECT 602.240 487.230 602.500 487.550 ;
        RECT 641.340 487.230 641.600 487.550 ;
        RECT 1376.480 19.370 1376.620 488.590 ;
        RECT 1376.420 19.050 1376.680 19.370 ;
        RECT 2024.100 18.710 2024.360 19.030 ;
        RECT 2024.160 2.400 2024.300 18.710 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
      LAYER via2 ;
        RECT 594.870 496.600 595.150 496.880 ;
        RECT 602.230 495.920 602.510 496.200 ;
      LAYER met3 ;
        RECT 594.845 496.890 595.175 496.905 ;
        RECT 594.845 496.590 602.290 496.890 ;
        RECT 594.845 496.575 595.175 496.590 ;
        RECT 601.990 496.225 602.290 496.590 ;
        RECT 601.990 495.910 602.535 496.225 ;
        RECT 602.205 495.895 602.535 495.910 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.390 116.180 594.710 116.240 ;
        RECT 2035.570 116.180 2035.890 116.240 ;
        RECT 594.390 116.040 2035.890 116.180 ;
        RECT 594.390 115.980 594.710 116.040 ;
        RECT 2035.570 115.980 2035.890 116.040 ;
        RECT 2035.570 16.900 2035.890 16.960 ;
        RECT 2042.010 16.900 2042.330 16.960 ;
        RECT 2035.570 16.760 2042.330 16.900 ;
        RECT 2035.570 16.700 2035.890 16.760 ;
        RECT 2042.010 16.700 2042.330 16.760 ;
      LAYER via ;
        RECT 594.420 115.980 594.680 116.240 ;
        RECT 2035.600 115.980 2035.860 116.240 ;
        RECT 2035.600 16.700 2035.860 16.960 ;
        RECT 2042.040 16.700 2042.300 16.960 ;
      LAYER met2 ;
        RECT 595.130 500.000 595.410 504.000 ;
        RECT 595.170 498.680 595.310 500.000 ;
        RECT 595.170 498.540 595.540 498.680 ;
        RECT 595.400 496.245 595.540 498.540 ;
        RECT 595.330 495.875 595.610 496.245 ;
        RECT 594.410 493.155 594.690 493.525 ;
        RECT 594.480 116.270 594.620 493.155 ;
        RECT 594.420 115.950 594.680 116.270 ;
        RECT 2035.600 115.950 2035.860 116.270 ;
        RECT 2035.660 16.990 2035.800 115.950 ;
        RECT 2035.600 16.670 2035.860 16.990 ;
        RECT 2042.040 16.670 2042.300 16.990 ;
        RECT 2042.100 2.400 2042.240 16.670 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
      LAYER via2 ;
        RECT 595.330 495.920 595.610 496.200 ;
        RECT 594.410 493.200 594.690 493.480 ;
      LAYER met3 ;
        RECT 594.590 496.210 594.970 496.220 ;
        RECT 595.305 496.210 595.635 496.225 ;
        RECT 594.590 495.910 595.635 496.210 ;
        RECT 594.590 495.900 594.970 495.910 ;
        RECT 595.305 495.895 595.635 495.910 ;
        RECT 594.385 493.500 594.715 493.505 ;
        RECT 594.385 493.490 594.970 493.500 ;
        RECT 594.160 493.190 594.970 493.490 ;
        RECT 594.385 493.180 594.970 493.190 ;
        RECT 594.385 493.175 594.715 493.180 ;
      LAYER via3 ;
        RECT 594.620 495.900 594.940 496.220 ;
        RECT 594.620 493.180 594.940 493.500 ;
      LAYER met4 ;
        RECT 594.615 495.895 594.945 496.225 ;
        RECT 594.630 493.505 594.930 495.895 ;
        RECT 594.615 493.175 594.945 493.505 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 495.720 499.160 496.040 499.420 ;
        RECT 495.030 497.660 495.350 497.720 ;
        RECT 495.810 497.660 495.950 499.160 ;
        RECT 495.030 497.520 495.950 497.660 ;
        RECT 495.030 497.460 495.350 497.520 ;
      LAYER via ;
        RECT 495.750 499.160 496.010 499.420 ;
        RECT 495.060 497.460 495.320 497.720 ;
      LAYER met2 ;
        RECT 495.770 500.000 496.050 504.000 ;
        RECT 495.810 499.450 495.950 500.000 ;
        RECT 495.750 499.130 496.010 499.450 ;
        RECT 495.060 497.430 495.320 497.750 ;
        RECT 495.120 488.085 495.260 497.430 ;
        RECT 495.050 487.715 495.330 488.085 ;
        RECT 759.550 113.715 759.830 114.085 ;
        RECT 759.620 82.870 759.760 113.715 ;
        RECT 759.620 82.730 765.280 82.870 ;
        RECT 765.140 2.400 765.280 82.730 ;
        RECT 764.930 -4.800 765.490 2.400 ;
      LAYER via2 ;
        RECT 495.050 487.760 495.330 488.040 ;
        RECT 759.550 113.760 759.830 114.040 ;
      LAYER met3 ;
        RECT 494.310 488.050 494.690 488.060 ;
        RECT 495.025 488.050 495.355 488.065 ;
        RECT 494.310 487.750 495.355 488.050 ;
        RECT 494.310 487.740 494.690 487.750 ;
        RECT 495.025 487.735 495.355 487.750 ;
        RECT 494.310 114.050 494.690 114.060 ;
        RECT 759.525 114.050 759.855 114.065 ;
        RECT 494.310 113.750 759.855 114.050 ;
        RECT 494.310 113.740 494.690 113.750 ;
        RECT 759.525 113.735 759.855 113.750 ;
      LAYER via3 ;
        RECT 494.340 487.740 494.660 488.060 ;
        RECT 494.340 113.740 494.660 114.060 ;
      LAYER met4 ;
        RECT 494.335 487.735 494.665 488.065 ;
        RECT 494.350 114.065 494.650 487.735 ;
        RECT 494.335 113.735 494.665 114.065 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 666.150 121.620 666.470 121.680 ;
        RECT 2056.270 121.620 2056.590 121.680 ;
        RECT 666.150 121.480 2056.590 121.620 ;
        RECT 666.150 121.420 666.470 121.480 ;
        RECT 2056.270 121.420 2056.590 121.480 ;
      LAYER via ;
        RECT 666.180 121.420 666.440 121.680 ;
        RECT 2056.300 121.420 2056.560 121.680 ;
      LAYER met2 ;
        RECT 596.510 500.000 596.790 504.000 ;
        RECT 596.550 499.815 596.690 500.000 ;
        RECT 596.480 499.445 596.760 499.815 ;
        RECT 598.090 497.915 598.370 498.285 ;
        RECT 598.160 488.765 598.300 497.915 ;
        RECT 598.090 488.395 598.370 488.765 ;
        RECT 665.710 488.395 665.990 488.765 ;
        RECT 665.780 487.290 665.920 488.395 ;
        RECT 665.780 487.150 666.380 487.290 ;
        RECT 666.240 121.710 666.380 487.150 ;
        RECT 666.180 121.390 666.440 121.710 ;
        RECT 2056.300 121.390 2056.560 121.710 ;
        RECT 2056.360 82.870 2056.500 121.390 ;
        RECT 2056.360 82.730 2059.720 82.870 ;
        RECT 2059.580 2.400 2059.720 82.730 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
      LAYER via2 ;
        RECT 596.480 499.490 596.760 499.770 ;
        RECT 598.090 497.960 598.370 498.240 ;
        RECT 598.090 488.440 598.370 488.720 ;
        RECT 665.710 488.440 665.990 488.720 ;
      LAYER met3 ;
        RECT 596.455 499.465 596.785 499.795 ;
        RECT 596.470 498.250 596.770 499.465 ;
        RECT 598.065 498.250 598.395 498.265 ;
        RECT 596.470 497.950 598.395 498.250 ;
        RECT 598.065 497.935 598.395 497.950 ;
        RECT 598.065 488.730 598.395 488.745 ;
        RECT 665.685 488.730 666.015 488.745 ;
        RECT 598.065 488.430 666.015 488.730 ;
        RECT 598.065 488.415 598.395 488.430 ;
        RECT 665.685 488.415 666.015 488.430 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 596.230 472.500 596.550 472.560 ;
        RECT 597.610 472.500 597.930 472.560 ;
        RECT 596.230 472.360 597.930 472.500 ;
        RECT 596.230 472.300 596.550 472.360 ;
        RECT 597.610 472.300 597.930 472.360 ;
        RECT 596.230 155.620 596.550 155.680 ;
        RECT 2076.970 155.620 2077.290 155.680 ;
        RECT 596.230 155.480 2077.290 155.620 ;
        RECT 596.230 155.420 596.550 155.480 ;
        RECT 2076.970 155.420 2077.290 155.480 ;
      LAYER via ;
        RECT 596.260 472.300 596.520 472.560 ;
        RECT 597.640 472.300 597.900 472.560 ;
        RECT 596.260 155.420 596.520 155.680 ;
        RECT 2077.000 155.420 2077.260 155.680 ;
      LAYER met2 ;
        RECT 597.890 500.000 598.170 504.000 ;
        RECT 597.930 498.680 598.070 500.000 ;
        RECT 597.700 498.540 598.070 498.680 ;
        RECT 597.700 472.590 597.840 498.540 ;
        RECT 596.260 472.270 596.520 472.590 ;
        RECT 597.640 472.270 597.900 472.590 ;
        RECT 596.320 155.710 596.460 472.270 ;
        RECT 596.260 155.390 596.520 155.710 ;
        RECT 2077.000 155.390 2077.260 155.710 ;
        RECT 2077.060 16.050 2077.200 155.390 ;
        RECT 2077.060 15.910 2077.660 16.050 ;
        RECT 2077.520 2.400 2077.660 15.910 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 667.070 176.360 667.390 176.420 ;
        RECT 2090.770 176.360 2091.090 176.420 ;
        RECT 667.070 176.220 2091.090 176.360 ;
        RECT 667.070 176.160 667.390 176.220 ;
        RECT 2090.770 176.160 2091.090 176.220 ;
      LAYER via ;
        RECT 667.100 176.160 667.360 176.420 ;
        RECT 2090.800 176.160 2091.060 176.420 ;
      LAYER met2 ;
        RECT 599.270 500.000 599.550 504.000 ;
        RECT 599.310 498.680 599.450 500.000 ;
        RECT 599.310 498.540 599.680 498.680 ;
        RECT 599.540 486.045 599.680 498.540 ;
        RECT 599.470 485.675 599.750 486.045 ;
        RECT 667.090 484.995 667.370 485.365 ;
        RECT 667.160 176.450 667.300 484.995 ;
        RECT 667.100 176.130 667.360 176.450 ;
        RECT 2090.800 176.130 2091.060 176.450 ;
        RECT 2090.860 82.870 2091.000 176.130 ;
        RECT 2090.860 82.730 2092.840 82.870 ;
        RECT 2092.700 1.770 2092.840 82.730 ;
        RECT 2094.790 1.770 2095.350 2.400 ;
        RECT 2092.700 1.630 2095.350 1.770 ;
        RECT 2094.790 -4.800 2095.350 1.630 ;
      LAYER via2 ;
        RECT 599.470 485.720 599.750 486.000 ;
        RECT 667.090 485.040 667.370 485.320 ;
      LAYER met3 ;
        RECT 599.445 486.010 599.775 486.025 ;
        RECT 599.445 485.710 661.170 486.010 ;
        RECT 599.445 485.695 599.775 485.710 ;
        RECT 660.870 485.330 661.170 485.710 ;
        RECT 667.065 485.330 667.395 485.345 ;
        RECT 660.870 485.030 667.395 485.330 ;
        RECT 667.065 485.015 667.395 485.030 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.600 499.500 600.920 499.760 ;
        RECT 600.690 499.020 600.830 499.500 ;
        RECT 600.690 498.880 601.520 499.020 ;
        RECT 601.380 498.400 601.520 498.880 ;
        RECT 601.290 498.140 601.610 498.400 ;
        RECT 602.670 169.900 602.990 169.960 ;
        RECT 2111.470 169.900 2111.790 169.960 ;
        RECT 602.670 169.760 2111.790 169.900 ;
        RECT 602.670 169.700 602.990 169.760 ;
        RECT 2111.470 169.700 2111.790 169.760 ;
      LAYER via ;
        RECT 600.630 499.500 600.890 499.760 ;
        RECT 601.320 498.140 601.580 498.400 ;
        RECT 602.700 169.700 602.960 169.960 ;
        RECT 2111.500 169.700 2111.760 169.960 ;
      LAYER met2 ;
        RECT 600.650 500.000 600.930 504.000 ;
        RECT 600.690 499.790 600.830 500.000 ;
        RECT 600.630 499.470 600.890 499.790 ;
        RECT 601.320 498.340 601.580 498.430 ;
        RECT 601.320 498.200 601.980 498.340 ;
        RECT 601.320 498.110 601.580 498.200 ;
        RECT 601.840 473.520 601.980 498.200 ;
        RECT 601.840 473.380 602.440 473.520 ;
        RECT 602.300 472.330 602.440 473.380 ;
        RECT 602.300 472.190 602.900 472.330 ;
        RECT 602.760 169.990 602.900 472.190 ;
        RECT 602.700 169.670 602.960 169.990 ;
        RECT 2111.500 169.670 2111.760 169.990 ;
        RECT 2111.560 82.870 2111.700 169.670 ;
        RECT 2111.560 82.730 2113.080 82.870 ;
        RECT 2112.940 2.400 2113.080 82.730 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 601.980 499.160 602.300 499.420 ;
        RECT 602.070 497.320 602.210 499.160 ;
        RECT 607.270 497.320 607.590 497.380 ;
        RECT 602.070 497.180 607.590 497.320 ;
        RECT 607.270 497.120 607.590 497.180 ;
        RECT 607.270 484.400 607.590 484.460 ;
        RECT 666.610 484.400 666.930 484.460 ;
        RECT 607.270 484.260 666.930 484.400 ;
        RECT 607.270 484.200 607.590 484.260 ;
        RECT 666.610 484.200 666.930 484.260 ;
        RECT 666.610 258.640 666.930 258.700 ;
        RECT 2125.270 258.640 2125.590 258.700 ;
        RECT 666.610 258.500 2125.590 258.640 ;
        RECT 666.610 258.440 666.930 258.500 ;
        RECT 2125.270 258.440 2125.590 258.500 ;
      LAYER via ;
        RECT 602.010 499.160 602.270 499.420 ;
        RECT 607.300 497.120 607.560 497.380 ;
        RECT 607.300 484.200 607.560 484.460 ;
        RECT 666.640 484.200 666.900 484.460 ;
        RECT 666.640 258.440 666.900 258.700 ;
        RECT 2125.300 258.440 2125.560 258.700 ;
      LAYER met2 ;
        RECT 602.030 500.000 602.310 504.000 ;
        RECT 602.070 499.450 602.210 500.000 ;
        RECT 602.010 499.130 602.270 499.450 ;
        RECT 607.300 497.090 607.560 497.410 ;
        RECT 607.360 484.490 607.500 497.090 ;
        RECT 607.300 484.170 607.560 484.490 ;
        RECT 666.640 484.170 666.900 484.490 ;
        RECT 666.700 258.730 666.840 484.170 ;
        RECT 666.640 258.410 666.900 258.730 ;
        RECT 2125.300 258.410 2125.560 258.730 ;
        RECT 2125.360 82.870 2125.500 258.410 ;
        RECT 2125.360 82.730 2128.720 82.870 ;
        RECT 2128.580 1.770 2128.720 82.730 ;
        RECT 2130.670 1.770 2131.230 2.400 ;
        RECT 2128.580 1.630 2131.230 1.770 ;
        RECT 2130.670 -4.800 2131.230 1.630 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 603.360 499.500 603.680 499.760 ;
        RECT 603.450 498.060 603.590 499.500 ;
        RECT 603.130 497.860 603.590 498.060 ;
        RECT 603.130 497.800 603.450 497.860 ;
        RECT 603.130 169.560 603.450 169.620 ;
        RECT 2145.970 169.560 2146.290 169.620 ;
        RECT 603.130 169.420 2146.290 169.560 ;
        RECT 603.130 169.360 603.450 169.420 ;
        RECT 2145.970 169.360 2146.290 169.420 ;
      LAYER via ;
        RECT 603.390 499.500 603.650 499.760 ;
        RECT 603.160 497.800 603.420 498.060 ;
        RECT 603.160 169.360 603.420 169.620 ;
        RECT 2146.000 169.360 2146.260 169.620 ;
      LAYER met2 ;
        RECT 603.410 500.000 603.690 504.000 ;
        RECT 603.450 499.790 603.590 500.000 ;
        RECT 603.390 499.470 603.650 499.790 ;
        RECT 603.160 497.770 603.420 498.090 ;
        RECT 603.220 169.650 603.360 497.770 ;
        RECT 603.160 169.330 603.420 169.650 ;
        RECT 2146.000 169.330 2146.260 169.650 ;
        RECT 2146.060 1.770 2146.200 169.330 ;
        RECT 2148.150 1.770 2148.710 2.400 ;
        RECT 2146.060 1.630 2148.710 1.770 ;
        RECT 2148.150 -4.800 2148.710 1.630 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 604.740 498.820 605.060 499.080 ;
        RECT 604.830 498.340 604.970 498.820 ;
        RECT 604.830 498.200 606.580 498.340 ;
        RECT 606.440 497.660 606.580 498.200 ;
        RECT 608.190 497.660 608.510 497.720 ;
        RECT 606.440 497.520 608.510 497.660 ;
        RECT 608.190 497.460 608.510 497.520 ;
        RECT 608.190 488.820 608.510 488.880 ;
        RECT 636.250 488.820 636.570 488.880 ;
        RECT 608.190 488.680 636.570 488.820 ;
        RECT 608.190 488.620 608.510 488.680 ;
        RECT 636.250 488.620 636.570 488.680 ;
        RECT 636.250 486.440 636.570 486.500 ;
        RECT 636.250 486.300 639.700 486.440 ;
        RECT 636.250 486.240 636.570 486.300 ;
        RECT 639.560 486.100 639.700 486.300 ;
        RECT 673.050 486.100 673.370 486.160 ;
        RECT 639.560 485.960 673.370 486.100 ;
        RECT 673.050 485.900 673.370 485.960 ;
        RECT 673.050 72.660 673.370 72.720 ;
        RECT 2160.230 72.660 2160.550 72.720 ;
        RECT 673.050 72.520 2160.550 72.660 ;
        RECT 673.050 72.460 673.370 72.520 ;
        RECT 2160.230 72.460 2160.550 72.520 ;
        RECT 2160.230 16.900 2160.550 16.960 ;
        RECT 2166.210 16.900 2166.530 16.960 ;
        RECT 2160.230 16.760 2166.530 16.900 ;
        RECT 2160.230 16.700 2160.550 16.760 ;
        RECT 2166.210 16.700 2166.530 16.760 ;
      LAYER via ;
        RECT 604.770 498.820 605.030 499.080 ;
        RECT 608.220 497.460 608.480 497.720 ;
        RECT 608.220 488.620 608.480 488.880 ;
        RECT 636.280 488.620 636.540 488.880 ;
        RECT 636.280 486.240 636.540 486.500 ;
        RECT 673.080 485.900 673.340 486.160 ;
        RECT 673.080 72.460 673.340 72.720 ;
        RECT 2160.260 72.460 2160.520 72.720 ;
        RECT 2160.260 16.700 2160.520 16.960 ;
        RECT 2166.240 16.700 2166.500 16.960 ;
      LAYER met2 ;
        RECT 604.790 500.000 605.070 504.000 ;
        RECT 604.830 499.110 604.970 500.000 ;
        RECT 604.770 498.790 605.030 499.110 ;
        RECT 608.220 497.430 608.480 497.750 ;
        RECT 608.280 488.910 608.420 497.430 ;
        RECT 608.220 488.590 608.480 488.910 ;
        RECT 636.280 488.590 636.540 488.910 ;
        RECT 636.340 486.530 636.480 488.590 ;
        RECT 636.280 486.210 636.540 486.530 ;
        RECT 673.080 485.870 673.340 486.190 ;
        RECT 673.140 72.750 673.280 485.870 ;
        RECT 673.080 72.430 673.340 72.750 ;
        RECT 2160.260 72.430 2160.520 72.750 ;
        RECT 2160.320 16.990 2160.460 72.430 ;
        RECT 2160.260 16.670 2160.520 16.990 ;
        RECT 2166.240 16.670 2166.500 16.990 ;
        RECT 2166.300 2.400 2166.440 16.670 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 606.120 499.500 606.440 499.760 ;
        RECT 606.210 499.080 606.350 499.500 ;
        RECT 605.890 498.880 606.350 499.080 ;
        RECT 605.890 498.820 606.210 498.880 ;
      LAYER via ;
        RECT 606.150 499.500 606.410 499.760 ;
        RECT 605.920 498.820 606.180 499.080 ;
      LAYER met2 ;
        RECT 606.170 500.000 606.450 504.000 ;
        RECT 606.210 499.790 606.350 500.000 ;
        RECT 606.150 499.470 606.410 499.790 ;
        RECT 605.920 498.790 606.180 499.110 ;
        RECT 605.980 498.170 606.120 498.790 ;
        RECT 605.520 498.030 606.120 498.170 ;
        RECT 605.520 498.000 605.660 498.030 ;
        RECT 605.060 497.860 605.660 498.000 ;
        RECT 605.060 488.085 605.200 497.860 ;
        RECT 604.990 487.715 605.270 488.085 ;
        RECT 2180.490 177.635 2180.770 178.005 ;
        RECT 2180.560 82.870 2180.700 177.635 ;
        RECT 2180.560 82.730 2183.920 82.870 ;
        RECT 2183.780 2.400 2183.920 82.730 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
      LAYER via2 ;
        RECT 604.990 487.760 605.270 488.040 ;
        RECT 2180.490 177.680 2180.770 177.960 ;
      LAYER met3 ;
        RECT 603.790 488.050 604.170 488.060 ;
        RECT 604.965 488.050 605.295 488.065 ;
        RECT 603.790 487.750 605.295 488.050 ;
        RECT 603.790 487.740 604.170 487.750 ;
        RECT 604.965 487.735 605.295 487.750 ;
        RECT 603.790 177.970 604.170 177.980 ;
        RECT 2180.465 177.970 2180.795 177.985 ;
        RECT 603.790 177.670 2180.795 177.970 ;
        RECT 603.790 177.660 604.170 177.670 ;
        RECT 2180.465 177.655 2180.795 177.670 ;
      LAYER via3 ;
        RECT 603.820 487.740 604.140 488.060 ;
        RECT 603.820 177.660 604.140 177.980 ;
      LAYER met4 ;
        RECT 603.815 487.735 604.145 488.065 ;
        RECT 603.830 177.985 604.130 487.735 ;
        RECT 603.815 177.655 604.145 177.985 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.500 499.700 607.820 499.760 ;
        RECT 607.500 499.560 610.950 499.700 ;
        RECT 607.500 499.500 607.820 499.560 ;
        RECT 610.810 496.980 610.950 499.560 ;
        RECT 626.130 497.320 626.450 497.380 ;
        RECT 625.300 497.180 626.450 497.320 ;
        RECT 625.300 496.980 625.440 497.180 ;
        RECT 626.130 497.120 626.450 497.180 ;
        RECT 610.810 496.840 625.440 496.980 ;
        RECT 626.130 485.760 626.450 485.820 ;
        RECT 636.250 485.760 636.570 485.820 ;
        RECT 626.130 485.620 636.570 485.760 ;
        RECT 626.130 485.560 626.450 485.620 ;
        RECT 636.250 485.560 636.570 485.620 ;
        RECT 636.250 485.080 636.570 485.140 ;
        RECT 673.970 485.080 674.290 485.140 ;
        RECT 636.250 484.940 674.290 485.080 ;
        RECT 636.250 484.880 636.570 484.940 ;
        RECT 673.970 484.880 674.290 484.940 ;
        RECT 673.970 182.820 674.290 182.880 ;
        RECT 2201.630 182.820 2201.950 182.880 ;
        RECT 673.970 182.680 2201.950 182.820 ;
        RECT 673.970 182.620 674.290 182.680 ;
        RECT 2201.630 182.620 2201.950 182.680 ;
      LAYER via ;
        RECT 607.530 499.500 607.790 499.760 ;
        RECT 626.160 497.120 626.420 497.380 ;
        RECT 626.160 485.560 626.420 485.820 ;
        RECT 636.280 485.560 636.540 485.820 ;
        RECT 636.280 484.880 636.540 485.140 ;
        RECT 674.000 484.880 674.260 485.140 ;
        RECT 674.000 182.620 674.260 182.880 ;
        RECT 2201.660 182.620 2201.920 182.880 ;
      LAYER met2 ;
        RECT 607.550 500.000 607.830 504.000 ;
        RECT 607.590 499.790 607.730 500.000 ;
        RECT 607.530 499.470 607.790 499.790 ;
        RECT 626.160 497.090 626.420 497.410 ;
        RECT 626.220 485.850 626.360 497.090 ;
        RECT 626.160 485.530 626.420 485.850 ;
        RECT 636.280 485.530 636.540 485.850 ;
        RECT 636.340 485.170 636.480 485.530 ;
        RECT 636.280 484.850 636.540 485.170 ;
        RECT 674.000 484.850 674.260 485.170 ;
        RECT 674.060 182.910 674.200 484.850 ;
        RECT 674.000 182.590 674.260 182.910 ;
        RECT 2201.660 182.590 2201.920 182.910 ;
        RECT 2201.720 2.400 2201.860 182.590 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 610.030 189.620 610.350 189.680 ;
        RECT 2214.970 189.620 2215.290 189.680 ;
        RECT 610.030 189.480 2215.290 189.620 ;
        RECT 610.030 189.420 610.350 189.480 ;
        RECT 2214.970 189.420 2215.290 189.480 ;
      LAYER via ;
        RECT 610.060 189.420 610.320 189.680 ;
        RECT 2215.000 189.420 2215.260 189.680 ;
      LAYER met2 ;
        RECT 608.930 500.000 609.210 504.000 ;
        RECT 608.970 499.645 609.110 500.000 ;
        RECT 608.900 499.275 609.180 499.645 ;
        RECT 610.510 497.915 610.790 498.285 ;
        RECT 610.580 420.970 610.720 497.915 ;
        RECT 610.120 420.830 610.720 420.970 ;
        RECT 610.120 189.710 610.260 420.830 ;
        RECT 610.060 189.390 610.320 189.710 ;
        RECT 2215.000 189.390 2215.260 189.710 ;
        RECT 2215.060 82.870 2215.200 189.390 ;
        RECT 2215.060 82.730 2217.040 82.870 ;
        RECT 2216.900 1.770 2217.040 82.730 ;
        RECT 2218.990 1.770 2219.550 2.400 ;
        RECT 2216.900 1.630 2219.550 1.770 ;
        RECT 2218.990 -4.800 2219.550 1.630 ;
      LAYER via2 ;
        RECT 608.900 499.320 609.180 499.600 ;
        RECT 610.510 497.960 610.790 498.240 ;
      LAYER met3 ;
        RECT 608.875 499.610 609.205 499.625 ;
        RECT 608.875 499.310 610.570 499.610 ;
        RECT 608.875 499.295 609.205 499.310 ;
        RECT 610.270 498.265 610.570 499.310 ;
        RECT 610.270 497.950 610.815 498.265 ;
        RECT 610.485 497.935 610.815 497.950 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.870 497.800 497.190 498.060 ;
        RECT 496.960 496.640 497.100 497.800 ;
        RECT 502.850 496.640 503.170 496.700 ;
        RECT 496.960 496.500 503.170 496.640 ;
        RECT 502.850 496.440 503.170 496.500 ;
        RECT 502.850 488.140 503.170 488.200 ;
        RECT 508.370 488.140 508.690 488.200 ;
        RECT 502.850 488.000 508.690 488.140 ;
        RECT 502.850 487.940 503.170 488.000 ;
        RECT 508.370 487.940 508.690 488.000 ;
        RECT 507.910 178.060 508.230 178.120 ;
        RECT 779.770 178.060 780.090 178.120 ;
        RECT 507.910 177.920 780.090 178.060 ;
        RECT 507.910 177.860 508.230 177.920 ;
        RECT 779.770 177.860 780.090 177.920 ;
      LAYER via ;
        RECT 496.900 497.800 497.160 498.060 ;
        RECT 502.880 496.440 503.140 496.700 ;
        RECT 502.880 487.940 503.140 488.200 ;
        RECT 508.400 487.940 508.660 488.200 ;
        RECT 507.940 177.860 508.200 178.120 ;
        RECT 779.800 177.860 780.060 178.120 ;
      LAYER met2 ;
        RECT 497.150 500.000 497.430 504.000 ;
        RECT 497.190 498.680 497.330 500.000 ;
        RECT 496.960 498.540 497.330 498.680 ;
        RECT 496.960 498.090 497.100 498.540 ;
        RECT 496.900 497.770 497.160 498.090 ;
        RECT 502.880 496.410 503.140 496.730 ;
        RECT 502.940 488.230 503.080 496.410 ;
        RECT 502.880 487.910 503.140 488.230 ;
        RECT 508.400 487.910 508.660 488.230 ;
        RECT 508.460 448.570 508.600 487.910 ;
        RECT 508.000 448.430 508.600 448.570 ;
        RECT 508.000 178.150 508.140 448.430 ;
        RECT 507.940 177.830 508.200 178.150 ;
        RECT 779.800 177.830 780.060 178.150 ;
        RECT 779.860 82.870 780.000 177.830 ;
        RECT 779.860 82.730 780.920 82.870 ;
        RECT 780.780 1.770 780.920 82.730 ;
        RECT 782.870 1.770 783.430 2.400 ;
        RECT 780.780 1.630 783.430 1.770 ;
        RECT 782.870 -4.800 783.430 1.630 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 610.030 488.140 610.350 488.200 ;
        RECT 616.470 488.140 616.790 488.200 ;
        RECT 610.030 488.000 616.790 488.140 ;
        RECT 610.030 487.940 610.350 488.000 ;
        RECT 616.470 487.940 616.790 488.000 ;
        RECT 616.470 485.420 616.790 485.480 ;
        RECT 616.470 485.280 636.020 485.420 ;
        RECT 616.470 485.220 616.790 485.280 ;
        RECT 635.880 484.740 636.020 485.280 ;
        RECT 673.510 484.740 673.830 484.800 ;
        RECT 635.880 484.600 673.830 484.740 ;
        RECT 673.510 484.540 673.830 484.600 ;
        RECT 673.510 80.140 673.830 80.200 ;
        RECT 2237.050 80.140 2237.370 80.200 ;
        RECT 673.510 80.000 2237.370 80.140 ;
        RECT 673.510 79.940 673.830 80.000 ;
        RECT 2237.050 79.940 2237.370 80.000 ;
      LAYER via ;
        RECT 610.060 487.940 610.320 488.200 ;
        RECT 616.500 487.940 616.760 488.200 ;
        RECT 616.500 485.220 616.760 485.480 ;
        RECT 673.540 484.540 673.800 484.800 ;
        RECT 673.540 79.940 673.800 80.200 ;
        RECT 2237.080 79.940 2237.340 80.200 ;
      LAYER met2 ;
        RECT 610.310 500.000 610.590 504.000 ;
        RECT 610.350 498.680 610.490 500.000 ;
        RECT 610.120 498.540 610.490 498.680 ;
        RECT 610.120 488.230 610.260 498.540 ;
        RECT 610.060 487.910 610.320 488.230 ;
        RECT 616.500 487.910 616.760 488.230 ;
        RECT 616.560 485.510 616.700 487.910 ;
        RECT 616.500 485.190 616.760 485.510 ;
        RECT 673.540 484.510 673.800 484.830 ;
        RECT 673.600 80.230 673.740 484.510 ;
        RECT 673.540 79.910 673.800 80.230 ;
        RECT 2237.080 79.910 2237.340 80.230 ;
        RECT 2237.140 2.400 2237.280 79.910 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.690 500.000 611.970 504.000 ;
        RECT 611.730 498.850 611.870 500.000 ;
        RECT 611.500 498.710 611.870 498.850 ;
        RECT 611.500 483.325 611.640 498.710 ;
        RECT 611.430 482.955 611.710 483.325 ;
        RECT 2249.490 189.195 2249.770 189.565 ;
        RECT 2249.560 82.870 2249.700 189.195 ;
        RECT 2249.560 82.730 2254.760 82.870 ;
        RECT 2254.620 2.400 2254.760 82.730 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
      LAYER via2 ;
        RECT 611.430 483.000 611.710 483.280 ;
        RECT 2249.490 189.240 2249.770 189.520 ;
      LAYER met3 ;
        RECT 610.230 483.290 610.610 483.300 ;
        RECT 611.405 483.290 611.735 483.305 ;
        RECT 610.230 482.990 611.735 483.290 ;
        RECT 610.230 482.980 610.610 482.990 ;
        RECT 611.405 482.975 611.735 482.990 ;
        RECT 610.230 189.530 610.610 189.540 ;
        RECT 2249.465 189.530 2249.795 189.545 ;
        RECT 610.230 189.230 2249.795 189.530 ;
        RECT 610.230 189.220 610.610 189.230 ;
        RECT 2249.465 189.215 2249.795 189.230 ;
      LAYER via3 ;
        RECT 610.260 482.980 610.580 483.300 ;
        RECT 610.260 189.220 610.580 189.540 ;
      LAYER met4 ;
        RECT 610.255 482.975 610.585 483.305 ;
        RECT 610.270 189.545 610.570 482.975 ;
        RECT 610.255 189.215 610.585 189.545 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.070 500.000 613.350 504.000 ;
        RECT 613.110 498.850 613.250 500.000 ;
        RECT 613.110 498.710 613.940 498.850 ;
        RECT 613.800 488.085 613.940 498.710 ;
        RECT 613.730 487.715 614.010 488.085 ;
        RECT 2270.190 487.715 2270.470 488.085 ;
        RECT 2270.260 1.770 2270.400 487.715 ;
        RECT 2272.350 1.770 2272.910 2.400 ;
        RECT 2270.260 1.630 2272.910 1.770 ;
        RECT 2272.350 -4.800 2272.910 1.630 ;
      LAYER via2 ;
        RECT 613.730 487.760 614.010 488.040 ;
        RECT 2270.190 487.760 2270.470 488.040 ;
      LAYER met3 ;
        RECT 613.705 488.050 614.035 488.065 ;
        RECT 2270.165 488.050 2270.495 488.065 ;
        RECT 613.705 487.750 2270.495 488.050 ;
        RECT 613.705 487.735 614.035 487.750 ;
        RECT 2270.165 487.735 2270.495 487.750 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 614.630 480.660 614.950 480.720 ;
        RECT 617.390 480.660 617.710 480.720 ;
        RECT 614.630 480.520 617.710 480.660 ;
        RECT 614.630 480.460 614.950 480.520 ;
        RECT 617.390 480.460 617.710 480.520 ;
        RECT 617.390 362.340 617.710 362.400 ;
        RECT 2283.970 362.340 2284.290 362.400 ;
        RECT 617.390 362.200 2284.290 362.340 ;
        RECT 617.390 362.140 617.710 362.200 ;
        RECT 2283.970 362.140 2284.290 362.200 ;
        RECT 2283.970 16.900 2284.290 16.960 ;
        RECT 2290.410 16.900 2290.730 16.960 ;
        RECT 2283.970 16.760 2290.730 16.900 ;
        RECT 2283.970 16.700 2284.290 16.760 ;
        RECT 2290.410 16.700 2290.730 16.760 ;
      LAYER via ;
        RECT 614.660 480.460 614.920 480.720 ;
        RECT 617.420 480.460 617.680 480.720 ;
        RECT 617.420 362.140 617.680 362.400 ;
        RECT 2284.000 362.140 2284.260 362.400 ;
        RECT 2284.000 16.700 2284.260 16.960 ;
        RECT 2290.440 16.700 2290.700 16.960 ;
      LAYER met2 ;
        RECT 614.450 500.000 614.730 504.000 ;
        RECT 614.490 498.680 614.630 500.000 ;
        RECT 614.490 498.540 614.860 498.680 ;
        RECT 614.720 480.750 614.860 498.540 ;
        RECT 614.660 480.430 614.920 480.750 ;
        RECT 617.420 480.430 617.680 480.750 ;
        RECT 617.480 362.430 617.620 480.430 ;
        RECT 617.420 362.110 617.680 362.430 ;
        RECT 2284.000 362.110 2284.260 362.430 ;
        RECT 2284.060 16.990 2284.200 362.110 ;
        RECT 2284.000 16.670 2284.260 16.990 ;
        RECT 2290.440 16.670 2290.700 16.990 ;
        RECT 2290.500 2.400 2290.640 16.670 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 667.070 487.460 667.390 487.520 ;
        RECT 2300.990 487.460 2301.310 487.520 ;
        RECT 667.070 487.320 2301.310 487.460 ;
        RECT 667.070 487.260 667.390 487.320 ;
        RECT 2300.990 487.260 2301.310 487.320 ;
        RECT 652.810 487.120 653.130 487.180 ;
        RECT 635.880 486.980 653.130 487.120 ;
        RECT 616.930 486.440 617.250 486.500 ;
        RECT 635.880 486.440 636.020 486.980 ;
        RECT 652.810 486.920 653.130 486.980 ;
        RECT 616.930 486.300 636.020 486.440 ;
        RECT 616.930 486.240 617.250 486.300 ;
        RECT 652.810 485.760 653.130 485.820 ;
        RECT 667.070 485.760 667.390 485.820 ;
        RECT 652.810 485.620 667.390 485.760 ;
        RECT 652.810 485.560 653.130 485.620 ;
        RECT 667.070 485.560 667.390 485.620 ;
        RECT 2300.990 14.860 2301.310 14.920 ;
        RECT 2307.890 14.860 2308.210 14.920 ;
        RECT 2300.990 14.720 2308.210 14.860 ;
        RECT 2300.990 14.660 2301.310 14.720 ;
        RECT 2307.890 14.660 2308.210 14.720 ;
      LAYER via ;
        RECT 667.100 487.260 667.360 487.520 ;
        RECT 2301.020 487.260 2301.280 487.520 ;
        RECT 616.960 486.240 617.220 486.500 ;
        RECT 652.840 486.920 653.100 487.180 ;
        RECT 652.840 485.560 653.100 485.820 ;
        RECT 667.100 485.560 667.360 485.820 ;
        RECT 2301.020 14.660 2301.280 14.920 ;
        RECT 2307.920 14.660 2308.180 14.920 ;
      LAYER met2 ;
        RECT 615.830 500.000 616.110 504.000 ;
        RECT 615.870 499.700 616.010 500.000 ;
        RECT 615.870 499.560 616.240 499.700 ;
        RECT 616.100 499.530 616.240 499.560 ;
        RECT 616.100 499.390 616.470 499.530 ;
        RECT 616.330 498.850 616.470 499.390 ;
        RECT 616.330 498.710 616.700 498.850 ;
        RECT 616.560 488.650 616.700 498.710 ;
        RECT 616.560 488.510 617.160 488.650 ;
        RECT 617.020 486.530 617.160 488.510 ;
        RECT 667.100 487.230 667.360 487.550 ;
        RECT 2301.020 487.230 2301.280 487.550 ;
        RECT 652.840 486.890 653.100 487.210 ;
        RECT 616.960 486.210 617.220 486.530 ;
        RECT 652.900 485.850 653.040 486.890 ;
        RECT 667.160 485.850 667.300 487.230 ;
        RECT 652.840 485.530 653.100 485.850 ;
        RECT 667.100 485.530 667.360 485.850 ;
        RECT 2301.080 14.950 2301.220 487.230 ;
        RECT 2301.020 14.630 2301.280 14.950 ;
        RECT 2307.920 14.630 2308.180 14.950 ;
        RECT 2307.980 2.400 2308.120 14.630 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 617.850 369.140 618.170 369.200 ;
        RECT 2325.370 369.140 2325.690 369.200 ;
        RECT 617.850 369.000 2325.690 369.140 ;
        RECT 617.850 368.940 618.170 369.000 ;
        RECT 2325.370 368.940 2325.690 369.000 ;
      LAYER via ;
        RECT 617.880 368.940 618.140 369.200 ;
        RECT 2325.400 368.940 2325.660 369.200 ;
      LAYER met2 ;
        RECT 617.210 500.000 617.490 504.000 ;
        RECT 617.250 498.680 617.390 500.000 ;
        RECT 617.250 498.540 617.620 498.680 ;
        RECT 617.480 498.340 617.620 498.540 ;
        RECT 617.480 498.200 618.080 498.340 ;
        RECT 617.940 369.230 618.080 498.200 ;
        RECT 617.880 368.910 618.140 369.230 ;
        RECT 2325.400 368.910 2325.660 369.230 ;
        RECT 2325.460 34.570 2325.600 368.910 ;
        RECT 2325.460 34.430 2326.060 34.570 ;
        RECT 2325.920 2.400 2326.060 34.430 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 618.540 499.160 618.860 499.420 ;
        RECT 618.630 497.660 618.770 499.160 ;
        RECT 619.230 497.660 619.550 497.720 ;
        RECT 618.630 497.520 619.550 497.660 ;
        RECT 619.230 497.460 619.550 497.520 ;
        RECT 672.590 18.600 672.910 18.660 ;
        RECT 2343.310 18.600 2343.630 18.660 ;
        RECT 672.590 18.460 2343.630 18.600 ;
        RECT 672.590 18.400 672.910 18.460 ;
        RECT 2343.310 18.400 2343.630 18.460 ;
      LAYER via ;
        RECT 618.570 499.160 618.830 499.420 ;
        RECT 619.260 497.460 619.520 497.720 ;
        RECT 672.620 18.400 672.880 18.660 ;
        RECT 2343.340 18.400 2343.600 18.660 ;
      LAYER met2 ;
        RECT 618.590 500.000 618.870 504.000 ;
        RECT 618.630 499.450 618.770 500.000 ;
        RECT 618.570 499.130 618.830 499.450 ;
        RECT 619.260 497.430 619.520 497.750 ;
        RECT 619.320 496.925 619.460 497.430 ;
        RECT 617.410 496.555 617.690 496.925 ;
        RECT 619.250 496.555 619.530 496.925 ;
        RECT 617.480 489.445 617.620 496.555 ;
        RECT 617.410 489.075 617.690 489.445 ;
        RECT 672.610 489.075 672.890 489.445 ;
        RECT 672.680 18.690 672.820 489.075 ;
        RECT 672.620 18.370 672.880 18.690 ;
        RECT 2343.340 18.370 2343.600 18.690 ;
        RECT 2343.400 2.400 2343.540 18.370 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
      LAYER via2 ;
        RECT 617.410 496.600 617.690 496.880 ;
        RECT 619.250 496.600 619.530 496.880 ;
        RECT 617.410 489.120 617.690 489.400 ;
        RECT 672.610 489.120 672.890 489.400 ;
      LAYER met3 ;
        RECT 617.385 496.890 617.715 496.905 ;
        RECT 619.225 496.890 619.555 496.905 ;
        RECT 617.385 496.590 619.555 496.890 ;
        RECT 617.385 496.575 617.715 496.590 ;
        RECT 619.225 496.575 619.555 496.590 ;
        RECT 617.385 489.410 617.715 489.425 ;
        RECT 672.585 489.410 672.915 489.425 ;
        RECT 617.385 489.110 672.915 489.410 ;
        RECT 617.385 489.095 617.715 489.110 ;
        RECT 672.585 489.095 672.915 489.110 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.970 500.000 620.250 504.000 ;
        RECT 620.010 498.680 620.150 500.000 ;
        RECT 620.010 498.540 620.380 498.680 ;
        RECT 620.240 483.325 620.380 498.540 ;
        RECT 620.170 482.955 620.450 483.325 ;
        RECT 2359.890 410.195 2360.170 410.565 ;
        RECT 2359.960 82.870 2360.100 410.195 ;
        RECT 2359.960 82.730 2361.480 82.870 ;
        RECT 2361.340 2.400 2361.480 82.730 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
      LAYER via2 ;
        RECT 620.170 483.000 620.450 483.280 ;
        RECT 2359.890 410.240 2360.170 410.520 ;
      LAYER met3 ;
        RECT 620.145 483.300 620.475 483.305 ;
        RECT 620.145 483.290 620.730 483.300 ;
        RECT 619.920 482.990 620.730 483.290 ;
        RECT 620.145 482.980 620.730 482.990 ;
        RECT 620.145 482.975 620.475 482.980 ;
        RECT 620.350 410.530 620.730 410.540 ;
        RECT 2359.865 410.530 2360.195 410.545 ;
        RECT 620.350 410.230 2360.195 410.530 ;
        RECT 620.350 410.220 620.730 410.230 ;
        RECT 2359.865 410.215 2360.195 410.230 ;
      LAYER via3 ;
        RECT 620.380 482.980 620.700 483.300 ;
        RECT 620.380 410.220 620.700 410.540 ;
      LAYER met4 ;
        RECT 620.375 482.975 620.705 483.305 ;
        RECT 620.390 410.545 620.690 482.975 ;
        RECT 620.375 410.215 620.705 410.545 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.300 499.500 621.620 499.760 ;
        RECT 621.390 498.000 621.530 499.500 ;
        RECT 621.990 498.000 622.310 498.060 ;
        RECT 621.390 497.860 622.310 498.000 ;
        RECT 621.990 497.800 622.310 497.860 ;
        RECT 621.990 488.480 622.310 488.540 ;
        RECT 632.570 488.480 632.890 488.540 ;
        RECT 621.990 488.340 632.890 488.480 ;
        RECT 621.990 488.280 622.310 488.340 ;
        RECT 632.570 488.280 632.890 488.340 ;
        RECT 632.570 483.720 632.890 483.780 ;
        RECT 1438.490 483.720 1438.810 483.780 ;
        RECT 632.570 483.580 1438.810 483.720 ;
        RECT 632.570 483.520 632.890 483.580 ;
        RECT 1438.490 483.520 1438.810 483.580 ;
        RECT 1438.490 67.220 1438.810 67.280 ;
        RECT 2378.730 67.220 2379.050 67.280 ;
        RECT 1438.490 67.080 2379.050 67.220 ;
        RECT 1438.490 67.020 1438.810 67.080 ;
        RECT 2378.730 67.020 2379.050 67.080 ;
      LAYER via ;
        RECT 621.330 499.500 621.590 499.760 ;
        RECT 622.020 497.800 622.280 498.060 ;
        RECT 622.020 488.280 622.280 488.540 ;
        RECT 632.600 488.280 632.860 488.540 ;
        RECT 632.600 483.520 632.860 483.780 ;
        RECT 1438.520 483.520 1438.780 483.780 ;
        RECT 1438.520 67.020 1438.780 67.280 ;
        RECT 2378.760 67.020 2379.020 67.280 ;
      LAYER met2 ;
        RECT 621.350 500.000 621.630 504.000 ;
        RECT 621.390 499.790 621.530 500.000 ;
        RECT 621.330 499.470 621.590 499.790 ;
        RECT 622.020 497.770 622.280 498.090 ;
        RECT 622.080 488.570 622.220 497.770 ;
        RECT 622.020 488.250 622.280 488.570 ;
        RECT 632.600 488.250 632.860 488.570 ;
        RECT 632.660 483.810 632.800 488.250 ;
        RECT 632.600 483.490 632.860 483.810 ;
        RECT 1438.520 483.490 1438.780 483.810 ;
        RECT 1438.580 67.310 1438.720 483.490 ;
        RECT 1438.520 66.990 1438.780 67.310 ;
        RECT 2378.760 66.990 2379.020 67.310 ;
        RECT 2378.820 2.400 2378.960 66.990 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.680 499.500 623.000 499.760 ;
        RECT 621.530 497.660 621.850 497.720 ;
        RECT 622.770 497.660 622.910 499.500 ;
        RECT 621.530 497.520 622.910 497.660 ;
        RECT 621.530 497.460 621.850 497.520 ;
        RECT 621.530 484.060 621.850 484.120 ;
        RECT 660.630 484.060 660.950 484.120 ;
        RECT 621.530 483.920 660.950 484.060 ;
        RECT 621.530 483.860 621.850 483.920 ;
        RECT 660.630 483.860 660.950 483.920 ;
        RECT 660.630 18.260 660.950 18.320 ;
        RECT 2396.670 18.260 2396.990 18.320 ;
        RECT 660.630 18.120 2396.990 18.260 ;
        RECT 660.630 18.060 660.950 18.120 ;
        RECT 2396.670 18.060 2396.990 18.120 ;
      LAYER via ;
        RECT 622.710 499.500 622.970 499.760 ;
        RECT 621.560 497.460 621.820 497.720 ;
        RECT 621.560 483.860 621.820 484.120 ;
        RECT 660.660 483.860 660.920 484.120 ;
        RECT 660.660 18.060 660.920 18.320 ;
        RECT 2396.700 18.060 2396.960 18.320 ;
      LAYER met2 ;
        RECT 622.730 500.000 623.010 504.000 ;
        RECT 622.770 499.790 622.910 500.000 ;
        RECT 622.710 499.470 622.970 499.790 ;
        RECT 621.560 497.430 621.820 497.750 ;
        RECT 621.620 484.150 621.760 497.430 ;
        RECT 621.560 483.830 621.820 484.150 ;
        RECT 660.660 483.830 660.920 484.150 ;
        RECT 660.720 18.350 660.860 483.830 ;
        RECT 660.660 18.030 660.920 18.350 ;
        RECT 2396.700 18.030 2396.960 18.350 ;
        RECT 2396.760 2.400 2396.900 18.030 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.870 24.040 497.190 24.100 ;
        RECT 641.770 24.040 642.090 24.100 ;
        RECT 496.870 23.900 642.090 24.040 ;
        RECT 496.870 23.840 497.190 23.900 ;
        RECT 641.770 23.840 642.090 23.900 ;
        RECT 641.770 19.620 642.090 19.680 ;
        RECT 800.470 19.620 800.790 19.680 ;
        RECT 641.770 19.480 800.790 19.620 ;
        RECT 641.770 19.420 642.090 19.480 ;
        RECT 800.470 19.420 800.790 19.480 ;
      LAYER via ;
        RECT 496.900 23.840 497.160 24.100 ;
        RECT 641.800 23.840 642.060 24.100 ;
        RECT 641.800 19.420 642.060 19.680 ;
        RECT 800.500 19.420 800.760 19.680 ;
      LAYER met2 ;
        RECT 498.530 500.000 498.810 504.000 ;
        RECT 498.570 498.680 498.710 500.000 ;
        RECT 498.570 498.540 498.940 498.680 ;
        RECT 498.800 498.285 498.940 498.540 ;
        RECT 498.730 497.915 499.010 498.285 ;
        RECT 496.890 497.235 497.170 497.605 ;
        RECT 496.960 24.130 497.100 497.235 ;
        RECT 496.900 23.810 497.160 24.130 ;
        RECT 641.800 23.810 642.060 24.130 ;
        RECT 641.860 19.710 642.000 23.810 ;
        RECT 641.800 19.390 642.060 19.710 ;
        RECT 800.500 19.390 800.760 19.710 ;
        RECT 800.560 2.400 800.700 19.390 ;
        RECT 800.350 -4.800 800.910 2.400 ;
      LAYER via2 ;
        RECT 498.730 497.960 499.010 498.240 ;
        RECT 496.890 497.280 497.170 497.560 ;
      LAYER met3 ;
        RECT 498.705 497.935 499.035 498.265 ;
        RECT 496.865 497.570 497.195 497.585 ;
        RECT 498.720 497.570 499.020 497.935 ;
        RECT 496.865 497.270 499.020 497.570 ;
        RECT 496.865 497.255 497.195 497.270 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 661.780 499.700 662.100 499.760 ;
        RECT 663.850 499.700 664.170 499.760 ;
        RECT 661.780 499.560 664.170 499.700 ;
        RECT 661.780 499.500 662.100 499.560 ;
        RECT 663.850 499.500 664.170 499.560 ;
        RECT 2328.590 65.860 2328.910 65.920 ;
        RECT 2905.430 65.860 2905.750 65.920 ;
        RECT 2328.590 65.720 2905.750 65.860 ;
        RECT 2328.590 65.660 2328.910 65.720 ;
        RECT 2905.430 65.660 2905.750 65.720 ;
      LAYER via ;
        RECT 661.810 499.500 662.070 499.760 ;
        RECT 663.880 499.500 664.140 499.760 ;
        RECT 2328.620 65.660 2328.880 65.920 ;
        RECT 2905.460 65.660 2905.720 65.920 ;
      LAYER met2 ;
        RECT 661.830 500.000 662.110 504.000 ;
        RECT 661.870 499.790 662.010 500.000 ;
        RECT 661.810 499.470 662.070 499.790 ;
        RECT 663.880 499.470 664.140 499.790 ;
        RECT 663.940 487.405 664.080 499.470 ;
        RECT 663.870 487.035 664.150 487.405 ;
        RECT 2328.610 487.035 2328.890 487.405 ;
        RECT 2328.680 65.950 2328.820 487.035 ;
        RECT 2328.620 65.630 2328.880 65.950 ;
        RECT 2905.460 65.630 2905.720 65.950 ;
        RECT 2905.520 16.730 2905.660 65.630 ;
        RECT 2905.060 16.590 2905.660 16.730 ;
        RECT 2905.060 2.400 2905.200 16.590 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 663.870 487.080 664.150 487.360 ;
        RECT 2328.610 487.080 2328.890 487.360 ;
      LAYER met3 ;
        RECT 663.845 487.370 664.175 487.385 ;
        RECT 2328.585 487.370 2328.915 487.385 ;
        RECT 663.845 487.070 2328.915 487.370 ;
        RECT 663.845 487.055 664.175 487.070 ;
        RECT 2328.585 487.055 2328.915 487.070 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 662.470 483.380 662.790 483.440 ;
        RECT 679.490 483.380 679.810 483.440 ;
        RECT 662.470 483.240 679.810 483.380 ;
        RECT 662.470 483.180 662.790 483.240 ;
        RECT 679.490 483.180 679.810 483.240 ;
        RECT 679.490 286.180 679.810 286.240 ;
        RECT 2904.970 286.180 2905.290 286.240 ;
        RECT 679.490 286.040 2905.290 286.180 ;
        RECT 679.490 285.980 679.810 286.040 ;
        RECT 2904.970 285.980 2905.290 286.040 ;
        RECT 2904.970 17.580 2905.290 17.640 ;
        RECT 2909.110 17.580 2909.430 17.640 ;
        RECT 2904.970 17.440 2909.430 17.580 ;
        RECT 2904.970 17.380 2905.290 17.440 ;
        RECT 2909.110 17.380 2909.430 17.440 ;
      LAYER via ;
        RECT 662.500 483.180 662.760 483.440 ;
        RECT 679.520 483.180 679.780 483.440 ;
        RECT 679.520 285.980 679.780 286.240 ;
        RECT 2905.000 285.980 2905.260 286.240 ;
        RECT 2905.000 17.380 2905.260 17.640 ;
        RECT 2909.140 17.380 2909.400 17.640 ;
      LAYER met2 ;
        RECT 662.290 500.000 662.570 504.000 ;
        RECT 662.330 499.530 662.470 500.000 ;
        RECT 662.330 499.390 662.700 499.530 ;
        RECT 662.560 483.470 662.700 499.390 ;
        RECT 662.500 483.150 662.760 483.470 ;
        RECT 679.520 483.150 679.780 483.470 ;
        RECT 679.580 286.270 679.720 483.150 ;
        RECT 679.520 285.950 679.780 286.270 ;
        RECT 2905.000 285.950 2905.260 286.270 ;
        RECT 2905.060 17.670 2905.200 285.950 ;
        RECT 2905.000 17.350 2905.260 17.670 ;
        RECT 2909.140 17.350 2909.400 17.670 ;
        RECT 2909.200 1.770 2909.340 17.350 ;
        RECT 2910.830 1.770 2911.390 2.400 ;
        RECT 2909.200 1.630 2911.390 1.770 ;
        RECT 2910.830 -4.800 2911.390 1.630 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 664.310 491.880 664.630 491.940 ;
        RECT 670.290 491.880 670.610 491.940 ;
        RECT 664.310 491.740 670.610 491.880 ;
        RECT 664.310 491.680 664.630 491.740 ;
        RECT 670.290 491.680 670.610 491.740 ;
        RECT 670.290 487.800 670.610 487.860 ;
        RECT 2114.690 487.800 2115.010 487.860 ;
        RECT 670.290 487.660 2115.010 487.800 ;
        RECT 670.290 487.600 670.610 487.660 ;
        RECT 2114.690 487.600 2115.010 487.660 ;
        RECT 2114.690 18.940 2115.010 19.000 ;
        RECT 2916.930 18.940 2917.250 19.000 ;
        RECT 2114.690 18.800 2917.250 18.940 ;
        RECT 2114.690 18.740 2115.010 18.800 ;
        RECT 2916.930 18.740 2917.250 18.800 ;
      LAYER via ;
        RECT 664.340 491.680 664.600 491.940 ;
        RECT 670.320 491.680 670.580 491.940 ;
        RECT 670.320 487.600 670.580 487.860 ;
        RECT 2114.720 487.600 2114.980 487.860 ;
        RECT 2114.720 18.740 2114.980 19.000 ;
        RECT 2916.960 18.740 2917.220 19.000 ;
      LAYER met2 ;
        RECT 662.750 500.210 663.030 504.000 ;
        RECT 662.750 500.070 664.540 500.210 ;
        RECT 662.750 500.000 663.030 500.070 ;
        RECT 664.400 491.970 664.540 500.070 ;
        RECT 664.340 491.650 664.600 491.970 ;
        RECT 670.320 491.650 670.580 491.970 ;
        RECT 670.380 487.890 670.520 491.650 ;
        RECT 670.320 487.570 670.580 487.890 ;
        RECT 2114.720 487.570 2114.980 487.890 ;
        RECT 2114.780 19.030 2114.920 487.570 ;
        RECT 2114.720 18.710 2114.980 19.030 ;
        RECT 2916.960 18.710 2917.220 19.030 ;
        RECT 2917.020 2.400 2917.160 18.710 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
        RECT 8.970 -38.270 12.070 3557.950 ;
        RECT 188.970 -38.270 192.070 3557.950 ;
        RECT 368.970 -38.270 372.070 3557.950 ;
        RECT 548.970 810.000 552.070 3557.950 ;
        RECT 421.040 510.640 422.640 788.560 ;
        RECT 574.640 510.640 576.240 788.560 ;
        RECT 548.970 -38.270 552.070 490.000 ;
        RECT 728.970 -38.270 732.070 3557.950 ;
        RECT 908.970 -38.270 912.070 3557.950 ;
        RECT 1088.970 -38.270 1092.070 3557.950 ;
        RECT 1268.970 -38.270 1272.070 3557.950 ;
        RECT 1448.970 -38.270 1452.070 3557.950 ;
        RECT 1628.970 -38.270 1632.070 3557.950 ;
        RECT 1808.970 -38.270 1812.070 3557.950 ;
        RECT 1988.970 -38.270 1992.070 3557.950 ;
        RECT 2168.970 -38.270 2172.070 3557.950 ;
        RECT 2348.970 -38.270 2352.070 3557.950 ;
        RECT 2528.970 -38.270 2532.070 3557.950 ;
        RECT 2708.970 -38.270 2712.070 3557.950 ;
        RECT 2888.970 -38.270 2892.070 3557.950 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
      LAYER via4 ;
        RECT -9.870 3523.010 -8.690 3524.190 ;
        RECT -8.270 3523.010 -7.090 3524.190 ;
        RECT -9.870 3521.410 -8.690 3522.590 ;
        RECT -8.270 3521.410 -7.090 3522.590 ;
        RECT -9.870 3436.090 -8.690 3437.270 ;
        RECT -8.270 3436.090 -7.090 3437.270 ;
        RECT -9.870 3434.490 -8.690 3435.670 ;
        RECT -8.270 3434.490 -7.090 3435.670 ;
        RECT -9.870 3256.090 -8.690 3257.270 ;
        RECT -8.270 3256.090 -7.090 3257.270 ;
        RECT -9.870 3254.490 -8.690 3255.670 ;
        RECT -8.270 3254.490 -7.090 3255.670 ;
        RECT -9.870 3076.090 -8.690 3077.270 ;
        RECT -8.270 3076.090 -7.090 3077.270 ;
        RECT -9.870 3074.490 -8.690 3075.670 ;
        RECT -8.270 3074.490 -7.090 3075.670 ;
        RECT -9.870 2896.090 -8.690 2897.270 ;
        RECT -8.270 2896.090 -7.090 2897.270 ;
        RECT -9.870 2894.490 -8.690 2895.670 ;
        RECT -8.270 2894.490 -7.090 2895.670 ;
        RECT -9.870 2716.090 -8.690 2717.270 ;
        RECT -8.270 2716.090 -7.090 2717.270 ;
        RECT -9.870 2714.490 -8.690 2715.670 ;
        RECT -8.270 2714.490 -7.090 2715.670 ;
        RECT -9.870 2536.090 -8.690 2537.270 ;
        RECT -8.270 2536.090 -7.090 2537.270 ;
        RECT -9.870 2534.490 -8.690 2535.670 ;
        RECT -8.270 2534.490 -7.090 2535.670 ;
        RECT -9.870 2356.090 -8.690 2357.270 ;
        RECT -8.270 2356.090 -7.090 2357.270 ;
        RECT -9.870 2354.490 -8.690 2355.670 ;
        RECT -8.270 2354.490 -7.090 2355.670 ;
        RECT -9.870 2176.090 -8.690 2177.270 ;
        RECT -8.270 2176.090 -7.090 2177.270 ;
        RECT -9.870 2174.490 -8.690 2175.670 ;
        RECT -8.270 2174.490 -7.090 2175.670 ;
        RECT -9.870 1996.090 -8.690 1997.270 ;
        RECT -8.270 1996.090 -7.090 1997.270 ;
        RECT -9.870 1994.490 -8.690 1995.670 ;
        RECT -8.270 1994.490 -7.090 1995.670 ;
        RECT -9.870 1816.090 -8.690 1817.270 ;
        RECT -8.270 1816.090 -7.090 1817.270 ;
        RECT -9.870 1814.490 -8.690 1815.670 ;
        RECT -8.270 1814.490 -7.090 1815.670 ;
        RECT -9.870 1636.090 -8.690 1637.270 ;
        RECT -8.270 1636.090 -7.090 1637.270 ;
        RECT -9.870 1634.490 -8.690 1635.670 ;
        RECT -8.270 1634.490 -7.090 1635.670 ;
        RECT -9.870 1456.090 -8.690 1457.270 ;
        RECT -8.270 1456.090 -7.090 1457.270 ;
        RECT -9.870 1454.490 -8.690 1455.670 ;
        RECT -8.270 1454.490 -7.090 1455.670 ;
        RECT -9.870 1276.090 -8.690 1277.270 ;
        RECT -8.270 1276.090 -7.090 1277.270 ;
        RECT -9.870 1274.490 -8.690 1275.670 ;
        RECT -8.270 1274.490 -7.090 1275.670 ;
        RECT -9.870 1096.090 -8.690 1097.270 ;
        RECT -8.270 1096.090 -7.090 1097.270 ;
        RECT -9.870 1094.490 -8.690 1095.670 ;
        RECT -8.270 1094.490 -7.090 1095.670 ;
        RECT -9.870 916.090 -8.690 917.270 ;
        RECT -8.270 916.090 -7.090 917.270 ;
        RECT -9.870 914.490 -8.690 915.670 ;
        RECT -8.270 914.490 -7.090 915.670 ;
        RECT -9.870 736.090 -8.690 737.270 ;
        RECT -8.270 736.090 -7.090 737.270 ;
        RECT -9.870 734.490 -8.690 735.670 ;
        RECT -8.270 734.490 -7.090 735.670 ;
        RECT -9.870 556.090 -8.690 557.270 ;
        RECT -8.270 556.090 -7.090 557.270 ;
        RECT -9.870 554.490 -8.690 555.670 ;
        RECT -8.270 554.490 -7.090 555.670 ;
        RECT -9.870 376.090 -8.690 377.270 ;
        RECT -8.270 376.090 -7.090 377.270 ;
        RECT -9.870 374.490 -8.690 375.670 ;
        RECT -8.270 374.490 -7.090 375.670 ;
        RECT -9.870 196.090 -8.690 197.270 ;
        RECT -8.270 196.090 -7.090 197.270 ;
        RECT -9.870 194.490 -8.690 195.670 ;
        RECT -8.270 194.490 -7.090 195.670 ;
        RECT -9.870 16.090 -8.690 17.270 ;
        RECT -8.270 16.090 -7.090 17.270 ;
        RECT -9.870 14.490 -8.690 15.670 ;
        RECT -8.270 14.490 -7.090 15.670 ;
        RECT -9.870 -2.910 -8.690 -1.730 ;
        RECT -8.270 -2.910 -7.090 -1.730 ;
        RECT -9.870 -4.510 -8.690 -3.330 ;
        RECT -8.270 -4.510 -7.090 -3.330 ;
        RECT 9.130 3523.010 10.310 3524.190 ;
        RECT 10.730 3523.010 11.910 3524.190 ;
        RECT 9.130 3521.410 10.310 3522.590 ;
        RECT 10.730 3521.410 11.910 3522.590 ;
        RECT 9.130 3436.090 10.310 3437.270 ;
        RECT 10.730 3436.090 11.910 3437.270 ;
        RECT 9.130 3434.490 10.310 3435.670 ;
        RECT 10.730 3434.490 11.910 3435.670 ;
        RECT 9.130 3256.090 10.310 3257.270 ;
        RECT 10.730 3256.090 11.910 3257.270 ;
        RECT 9.130 3254.490 10.310 3255.670 ;
        RECT 10.730 3254.490 11.910 3255.670 ;
        RECT 9.130 3076.090 10.310 3077.270 ;
        RECT 10.730 3076.090 11.910 3077.270 ;
        RECT 9.130 3074.490 10.310 3075.670 ;
        RECT 10.730 3074.490 11.910 3075.670 ;
        RECT 9.130 2896.090 10.310 2897.270 ;
        RECT 10.730 2896.090 11.910 2897.270 ;
        RECT 9.130 2894.490 10.310 2895.670 ;
        RECT 10.730 2894.490 11.910 2895.670 ;
        RECT 9.130 2716.090 10.310 2717.270 ;
        RECT 10.730 2716.090 11.910 2717.270 ;
        RECT 9.130 2714.490 10.310 2715.670 ;
        RECT 10.730 2714.490 11.910 2715.670 ;
        RECT 9.130 2536.090 10.310 2537.270 ;
        RECT 10.730 2536.090 11.910 2537.270 ;
        RECT 9.130 2534.490 10.310 2535.670 ;
        RECT 10.730 2534.490 11.910 2535.670 ;
        RECT 9.130 2356.090 10.310 2357.270 ;
        RECT 10.730 2356.090 11.910 2357.270 ;
        RECT 9.130 2354.490 10.310 2355.670 ;
        RECT 10.730 2354.490 11.910 2355.670 ;
        RECT 9.130 2176.090 10.310 2177.270 ;
        RECT 10.730 2176.090 11.910 2177.270 ;
        RECT 9.130 2174.490 10.310 2175.670 ;
        RECT 10.730 2174.490 11.910 2175.670 ;
        RECT 9.130 1996.090 10.310 1997.270 ;
        RECT 10.730 1996.090 11.910 1997.270 ;
        RECT 9.130 1994.490 10.310 1995.670 ;
        RECT 10.730 1994.490 11.910 1995.670 ;
        RECT 9.130 1816.090 10.310 1817.270 ;
        RECT 10.730 1816.090 11.910 1817.270 ;
        RECT 9.130 1814.490 10.310 1815.670 ;
        RECT 10.730 1814.490 11.910 1815.670 ;
        RECT 9.130 1636.090 10.310 1637.270 ;
        RECT 10.730 1636.090 11.910 1637.270 ;
        RECT 9.130 1634.490 10.310 1635.670 ;
        RECT 10.730 1634.490 11.910 1635.670 ;
        RECT 9.130 1456.090 10.310 1457.270 ;
        RECT 10.730 1456.090 11.910 1457.270 ;
        RECT 9.130 1454.490 10.310 1455.670 ;
        RECT 10.730 1454.490 11.910 1455.670 ;
        RECT 9.130 1276.090 10.310 1277.270 ;
        RECT 10.730 1276.090 11.910 1277.270 ;
        RECT 9.130 1274.490 10.310 1275.670 ;
        RECT 10.730 1274.490 11.910 1275.670 ;
        RECT 9.130 1096.090 10.310 1097.270 ;
        RECT 10.730 1096.090 11.910 1097.270 ;
        RECT 9.130 1094.490 10.310 1095.670 ;
        RECT 10.730 1094.490 11.910 1095.670 ;
        RECT 9.130 916.090 10.310 917.270 ;
        RECT 10.730 916.090 11.910 917.270 ;
        RECT 9.130 914.490 10.310 915.670 ;
        RECT 10.730 914.490 11.910 915.670 ;
        RECT 9.130 736.090 10.310 737.270 ;
        RECT 10.730 736.090 11.910 737.270 ;
        RECT 9.130 734.490 10.310 735.670 ;
        RECT 10.730 734.490 11.910 735.670 ;
        RECT 9.130 556.090 10.310 557.270 ;
        RECT 10.730 556.090 11.910 557.270 ;
        RECT 9.130 554.490 10.310 555.670 ;
        RECT 10.730 554.490 11.910 555.670 ;
        RECT 9.130 376.090 10.310 377.270 ;
        RECT 10.730 376.090 11.910 377.270 ;
        RECT 9.130 374.490 10.310 375.670 ;
        RECT 10.730 374.490 11.910 375.670 ;
        RECT 9.130 196.090 10.310 197.270 ;
        RECT 10.730 196.090 11.910 197.270 ;
        RECT 9.130 194.490 10.310 195.670 ;
        RECT 10.730 194.490 11.910 195.670 ;
        RECT 9.130 16.090 10.310 17.270 ;
        RECT 10.730 16.090 11.910 17.270 ;
        RECT 9.130 14.490 10.310 15.670 ;
        RECT 10.730 14.490 11.910 15.670 ;
        RECT 9.130 -2.910 10.310 -1.730 ;
        RECT 10.730 -2.910 11.910 -1.730 ;
        RECT 9.130 -4.510 10.310 -3.330 ;
        RECT 10.730 -4.510 11.910 -3.330 ;
        RECT 189.130 3523.010 190.310 3524.190 ;
        RECT 190.730 3523.010 191.910 3524.190 ;
        RECT 189.130 3521.410 190.310 3522.590 ;
        RECT 190.730 3521.410 191.910 3522.590 ;
        RECT 189.130 3436.090 190.310 3437.270 ;
        RECT 190.730 3436.090 191.910 3437.270 ;
        RECT 189.130 3434.490 190.310 3435.670 ;
        RECT 190.730 3434.490 191.910 3435.670 ;
        RECT 189.130 3256.090 190.310 3257.270 ;
        RECT 190.730 3256.090 191.910 3257.270 ;
        RECT 189.130 3254.490 190.310 3255.670 ;
        RECT 190.730 3254.490 191.910 3255.670 ;
        RECT 189.130 3076.090 190.310 3077.270 ;
        RECT 190.730 3076.090 191.910 3077.270 ;
        RECT 189.130 3074.490 190.310 3075.670 ;
        RECT 190.730 3074.490 191.910 3075.670 ;
        RECT 189.130 2896.090 190.310 2897.270 ;
        RECT 190.730 2896.090 191.910 2897.270 ;
        RECT 189.130 2894.490 190.310 2895.670 ;
        RECT 190.730 2894.490 191.910 2895.670 ;
        RECT 189.130 2716.090 190.310 2717.270 ;
        RECT 190.730 2716.090 191.910 2717.270 ;
        RECT 189.130 2714.490 190.310 2715.670 ;
        RECT 190.730 2714.490 191.910 2715.670 ;
        RECT 189.130 2536.090 190.310 2537.270 ;
        RECT 190.730 2536.090 191.910 2537.270 ;
        RECT 189.130 2534.490 190.310 2535.670 ;
        RECT 190.730 2534.490 191.910 2535.670 ;
        RECT 189.130 2356.090 190.310 2357.270 ;
        RECT 190.730 2356.090 191.910 2357.270 ;
        RECT 189.130 2354.490 190.310 2355.670 ;
        RECT 190.730 2354.490 191.910 2355.670 ;
        RECT 189.130 2176.090 190.310 2177.270 ;
        RECT 190.730 2176.090 191.910 2177.270 ;
        RECT 189.130 2174.490 190.310 2175.670 ;
        RECT 190.730 2174.490 191.910 2175.670 ;
        RECT 189.130 1996.090 190.310 1997.270 ;
        RECT 190.730 1996.090 191.910 1997.270 ;
        RECT 189.130 1994.490 190.310 1995.670 ;
        RECT 190.730 1994.490 191.910 1995.670 ;
        RECT 189.130 1816.090 190.310 1817.270 ;
        RECT 190.730 1816.090 191.910 1817.270 ;
        RECT 189.130 1814.490 190.310 1815.670 ;
        RECT 190.730 1814.490 191.910 1815.670 ;
        RECT 189.130 1636.090 190.310 1637.270 ;
        RECT 190.730 1636.090 191.910 1637.270 ;
        RECT 189.130 1634.490 190.310 1635.670 ;
        RECT 190.730 1634.490 191.910 1635.670 ;
        RECT 189.130 1456.090 190.310 1457.270 ;
        RECT 190.730 1456.090 191.910 1457.270 ;
        RECT 189.130 1454.490 190.310 1455.670 ;
        RECT 190.730 1454.490 191.910 1455.670 ;
        RECT 189.130 1276.090 190.310 1277.270 ;
        RECT 190.730 1276.090 191.910 1277.270 ;
        RECT 189.130 1274.490 190.310 1275.670 ;
        RECT 190.730 1274.490 191.910 1275.670 ;
        RECT 189.130 1096.090 190.310 1097.270 ;
        RECT 190.730 1096.090 191.910 1097.270 ;
        RECT 189.130 1094.490 190.310 1095.670 ;
        RECT 190.730 1094.490 191.910 1095.670 ;
        RECT 189.130 916.090 190.310 917.270 ;
        RECT 190.730 916.090 191.910 917.270 ;
        RECT 189.130 914.490 190.310 915.670 ;
        RECT 190.730 914.490 191.910 915.670 ;
        RECT 189.130 736.090 190.310 737.270 ;
        RECT 190.730 736.090 191.910 737.270 ;
        RECT 189.130 734.490 190.310 735.670 ;
        RECT 190.730 734.490 191.910 735.670 ;
        RECT 189.130 556.090 190.310 557.270 ;
        RECT 190.730 556.090 191.910 557.270 ;
        RECT 189.130 554.490 190.310 555.670 ;
        RECT 190.730 554.490 191.910 555.670 ;
        RECT 189.130 376.090 190.310 377.270 ;
        RECT 190.730 376.090 191.910 377.270 ;
        RECT 189.130 374.490 190.310 375.670 ;
        RECT 190.730 374.490 191.910 375.670 ;
        RECT 189.130 196.090 190.310 197.270 ;
        RECT 190.730 196.090 191.910 197.270 ;
        RECT 189.130 194.490 190.310 195.670 ;
        RECT 190.730 194.490 191.910 195.670 ;
        RECT 189.130 16.090 190.310 17.270 ;
        RECT 190.730 16.090 191.910 17.270 ;
        RECT 189.130 14.490 190.310 15.670 ;
        RECT 190.730 14.490 191.910 15.670 ;
        RECT 189.130 -2.910 190.310 -1.730 ;
        RECT 190.730 -2.910 191.910 -1.730 ;
        RECT 189.130 -4.510 190.310 -3.330 ;
        RECT 190.730 -4.510 191.910 -3.330 ;
        RECT 369.130 3523.010 370.310 3524.190 ;
        RECT 370.730 3523.010 371.910 3524.190 ;
        RECT 369.130 3521.410 370.310 3522.590 ;
        RECT 370.730 3521.410 371.910 3522.590 ;
        RECT 369.130 3436.090 370.310 3437.270 ;
        RECT 370.730 3436.090 371.910 3437.270 ;
        RECT 369.130 3434.490 370.310 3435.670 ;
        RECT 370.730 3434.490 371.910 3435.670 ;
        RECT 369.130 3256.090 370.310 3257.270 ;
        RECT 370.730 3256.090 371.910 3257.270 ;
        RECT 369.130 3254.490 370.310 3255.670 ;
        RECT 370.730 3254.490 371.910 3255.670 ;
        RECT 369.130 3076.090 370.310 3077.270 ;
        RECT 370.730 3076.090 371.910 3077.270 ;
        RECT 369.130 3074.490 370.310 3075.670 ;
        RECT 370.730 3074.490 371.910 3075.670 ;
        RECT 369.130 2896.090 370.310 2897.270 ;
        RECT 370.730 2896.090 371.910 2897.270 ;
        RECT 369.130 2894.490 370.310 2895.670 ;
        RECT 370.730 2894.490 371.910 2895.670 ;
        RECT 369.130 2716.090 370.310 2717.270 ;
        RECT 370.730 2716.090 371.910 2717.270 ;
        RECT 369.130 2714.490 370.310 2715.670 ;
        RECT 370.730 2714.490 371.910 2715.670 ;
        RECT 369.130 2536.090 370.310 2537.270 ;
        RECT 370.730 2536.090 371.910 2537.270 ;
        RECT 369.130 2534.490 370.310 2535.670 ;
        RECT 370.730 2534.490 371.910 2535.670 ;
        RECT 369.130 2356.090 370.310 2357.270 ;
        RECT 370.730 2356.090 371.910 2357.270 ;
        RECT 369.130 2354.490 370.310 2355.670 ;
        RECT 370.730 2354.490 371.910 2355.670 ;
        RECT 369.130 2176.090 370.310 2177.270 ;
        RECT 370.730 2176.090 371.910 2177.270 ;
        RECT 369.130 2174.490 370.310 2175.670 ;
        RECT 370.730 2174.490 371.910 2175.670 ;
        RECT 369.130 1996.090 370.310 1997.270 ;
        RECT 370.730 1996.090 371.910 1997.270 ;
        RECT 369.130 1994.490 370.310 1995.670 ;
        RECT 370.730 1994.490 371.910 1995.670 ;
        RECT 369.130 1816.090 370.310 1817.270 ;
        RECT 370.730 1816.090 371.910 1817.270 ;
        RECT 369.130 1814.490 370.310 1815.670 ;
        RECT 370.730 1814.490 371.910 1815.670 ;
        RECT 369.130 1636.090 370.310 1637.270 ;
        RECT 370.730 1636.090 371.910 1637.270 ;
        RECT 369.130 1634.490 370.310 1635.670 ;
        RECT 370.730 1634.490 371.910 1635.670 ;
        RECT 369.130 1456.090 370.310 1457.270 ;
        RECT 370.730 1456.090 371.910 1457.270 ;
        RECT 369.130 1454.490 370.310 1455.670 ;
        RECT 370.730 1454.490 371.910 1455.670 ;
        RECT 369.130 1276.090 370.310 1277.270 ;
        RECT 370.730 1276.090 371.910 1277.270 ;
        RECT 369.130 1274.490 370.310 1275.670 ;
        RECT 370.730 1274.490 371.910 1275.670 ;
        RECT 369.130 1096.090 370.310 1097.270 ;
        RECT 370.730 1096.090 371.910 1097.270 ;
        RECT 369.130 1094.490 370.310 1095.670 ;
        RECT 370.730 1094.490 371.910 1095.670 ;
        RECT 369.130 916.090 370.310 917.270 ;
        RECT 370.730 916.090 371.910 917.270 ;
        RECT 369.130 914.490 370.310 915.670 ;
        RECT 370.730 914.490 371.910 915.670 ;
        RECT 549.130 3523.010 550.310 3524.190 ;
        RECT 550.730 3523.010 551.910 3524.190 ;
        RECT 549.130 3521.410 550.310 3522.590 ;
        RECT 550.730 3521.410 551.910 3522.590 ;
        RECT 549.130 3436.090 550.310 3437.270 ;
        RECT 550.730 3436.090 551.910 3437.270 ;
        RECT 549.130 3434.490 550.310 3435.670 ;
        RECT 550.730 3434.490 551.910 3435.670 ;
        RECT 549.130 3256.090 550.310 3257.270 ;
        RECT 550.730 3256.090 551.910 3257.270 ;
        RECT 549.130 3254.490 550.310 3255.670 ;
        RECT 550.730 3254.490 551.910 3255.670 ;
        RECT 549.130 3076.090 550.310 3077.270 ;
        RECT 550.730 3076.090 551.910 3077.270 ;
        RECT 549.130 3074.490 550.310 3075.670 ;
        RECT 550.730 3074.490 551.910 3075.670 ;
        RECT 549.130 2896.090 550.310 2897.270 ;
        RECT 550.730 2896.090 551.910 2897.270 ;
        RECT 549.130 2894.490 550.310 2895.670 ;
        RECT 550.730 2894.490 551.910 2895.670 ;
        RECT 549.130 2716.090 550.310 2717.270 ;
        RECT 550.730 2716.090 551.910 2717.270 ;
        RECT 549.130 2714.490 550.310 2715.670 ;
        RECT 550.730 2714.490 551.910 2715.670 ;
        RECT 549.130 2536.090 550.310 2537.270 ;
        RECT 550.730 2536.090 551.910 2537.270 ;
        RECT 549.130 2534.490 550.310 2535.670 ;
        RECT 550.730 2534.490 551.910 2535.670 ;
        RECT 549.130 2356.090 550.310 2357.270 ;
        RECT 550.730 2356.090 551.910 2357.270 ;
        RECT 549.130 2354.490 550.310 2355.670 ;
        RECT 550.730 2354.490 551.910 2355.670 ;
        RECT 549.130 2176.090 550.310 2177.270 ;
        RECT 550.730 2176.090 551.910 2177.270 ;
        RECT 549.130 2174.490 550.310 2175.670 ;
        RECT 550.730 2174.490 551.910 2175.670 ;
        RECT 549.130 1996.090 550.310 1997.270 ;
        RECT 550.730 1996.090 551.910 1997.270 ;
        RECT 549.130 1994.490 550.310 1995.670 ;
        RECT 550.730 1994.490 551.910 1995.670 ;
        RECT 549.130 1816.090 550.310 1817.270 ;
        RECT 550.730 1816.090 551.910 1817.270 ;
        RECT 549.130 1814.490 550.310 1815.670 ;
        RECT 550.730 1814.490 551.910 1815.670 ;
        RECT 549.130 1636.090 550.310 1637.270 ;
        RECT 550.730 1636.090 551.910 1637.270 ;
        RECT 549.130 1634.490 550.310 1635.670 ;
        RECT 550.730 1634.490 551.910 1635.670 ;
        RECT 549.130 1456.090 550.310 1457.270 ;
        RECT 550.730 1456.090 551.910 1457.270 ;
        RECT 549.130 1454.490 550.310 1455.670 ;
        RECT 550.730 1454.490 551.910 1455.670 ;
        RECT 549.130 1276.090 550.310 1277.270 ;
        RECT 550.730 1276.090 551.910 1277.270 ;
        RECT 549.130 1274.490 550.310 1275.670 ;
        RECT 550.730 1274.490 551.910 1275.670 ;
        RECT 549.130 1096.090 550.310 1097.270 ;
        RECT 550.730 1096.090 551.910 1097.270 ;
        RECT 549.130 1094.490 550.310 1095.670 ;
        RECT 550.730 1094.490 551.910 1095.670 ;
        RECT 549.130 916.090 550.310 917.270 ;
        RECT 550.730 916.090 551.910 917.270 ;
        RECT 549.130 914.490 550.310 915.670 ;
        RECT 550.730 914.490 551.910 915.670 ;
        RECT 729.130 3523.010 730.310 3524.190 ;
        RECT 730.730 3523.010 731.910 3524.190 ;
        RECT 729.130 3521.410 730.310 3522.590 ;
        RECT 730.730 3521.410 731.910 3522.590 ;
        RECT 729.130 3436.090 730.310 3437.270 ;
        RECT 730.730 3436.090 731.910 3437.270 ;
        RECT 729.130 3434.490 730.310 3435.670 ;
        RECT 730.730 3434.490 731.910 3435.670 ;
        RECT 729.130 3256.090 730.310 3257.270 ;
        RECT 730.730 3256.090 731.910 3257.270 ;
        RECT 729.130 3254.490 730.310 3255.670 ;
        RECT 730.730 3254.490 731.910 3255.670 ;
        RECT 729.130 3076.090 730.310 3077.270 ;
        RECT 730.730 3076.090 731.910 3077.270 ;
        RECT 729.130 3074.490 730.310 3075.670 ;
        RECT 730.730 3074.490 731.910 3075.670 ;
        RECT 729.130 2896.090 730.310 2897.270 ;
        RECT 730.730 2896.090 731.910 2897.270 ;
        RECT 729.130 2894.490 730.310 2895.670 ;
        RECT 730.730 2894.490 731.910 2895.670 ;
        RECT 729.130 2716.090 730.310 2717.270 ;
        RECT 730.730 2716.090 731.910 2717.270 ;
        RECT 729.130 2714.490 730.310 2715.670 ;
        RECT 730.730 2714.490 731.910 2715.670 ;
        RECT 729.130 2536.090 730.310 2537.270 ;
        RECT 730.730 2536.090 731.910 2537.270 ;
        RECT 729.130 2534.490 730.310 2535.670 ;
        RECT 730.730 2534.490 731.910 2535.670 ;
        RECT 729.130 2356.090 730.310 2357.270 ;
        RECT 730.730 2356.090 731.910 2357.270 ;
        RECT 729.130 2354.490 730.310 2355.670 ;
        RECT 730.730 2354.490 731.910 2355.670 ;
        RECT 729.130 2176.090 730.310 2177.270 ;
        RECT 730.730 2176.090 731.910 2177.270 ;
        RECT 729.130 2174.490 730.310 2175.670 ;
        RECT 730.730 2174.490 731.910 2175.670 ;
        RECT 729.130 1996.090 730.310 1997.270 ;
        RECT 730.730 1996.090 731.910 1997.270 ;
        RECT 729.130 1994.490 730.310 1995.670 ;
        RECT 730.730 1994.490 731.910 1995.670 ;
        RECT 729.130 1816.090 730.310 1817.270 ;
        RECT 730.730 1816.090 731.910 1817.270 ;
        RECT 729.130 1814.490 730.310 1815.670 ;
        RECT 730.730 1814.490 731.910 1815.670 ;
        RECT 729.130 1636.090 730.310 1637.270 ;
        RECT 730.730 1636.090 731.910 1637.270 ;
        RECT 729.130 1634.490 730.310 1635.670 ;
        RECT 730.730 1634.490 731.910 1635.670 ;
        RECT 729.130 1456.090 730.310 1457.270 ;
        RECT 730.730 1456.090 731.910 1457.270 ;
        RECT 729.130 1454.490 730.310 1455.670 ;
        RECT 730.730 1454.490 731.910 1455.670 ;
        RECT 729.130 1276.090 730.310 1277.270 ;
        RECT 730.730 1276.090 731.910 1277.270 ;
        RECT 729.130 1274.490 730.310 1275.670 ;
        RECT 730.730 1274.490 731.910 1275.670 ;
        RECT 729.130 1096.090 730.310 1097.270 ;
        RECT 730.730 1096.090 731.910 1097.270 ;
        RECT 729.130 1094.490 730.310 1095.670 ;
        RECT 730.730 1094.490 731.910 1095.670 ;
        RECT 729.130 916.090 730.310 917.270 ;
        RECT 730.730 916.090 731.910 917.270 ;
        RECT 729.130 914.490 730.310 915.670 ;
        RECT 730.730 914.490 731.910 915.670 ;
        RECT 369.130 736.090 370.310 737.270 ;
        RECT 370.730 736.090 371.910 737.270 ;
        RECT 369.130 734.490 370.310 735.670 ;
        RECT 370.730 734.490 371.910 735.670 ;
        RECT 369.130 556.090 370.310 557.270 ;
        RECT 370.730 556.090 371.910 557.270 ;
        RECT 369.130 554.490 370.310 555.670 ;
        RECT 370.730 554.490 371.910 555.670 ;
        RECT 421.250 736.090 422.430 737.270 ;
        RECT 421.250 734.490 422.430 735.670 ;
        RECT 421.250 556.090 422.430 557.270 ;
        RECT 421.250 554.490 422.430 555.670 ;
        RECT 574.850 736.090 576.030 737.270 ;
        RECT 574.850 734.490 576.030 735.670 ;
        RECT 574.850 556.090 576.030 557.270 ;
        RECT 574.850 554.490 576.030 555.670 ;
        RECT 729.130 736.090 730.310 737.270 ;
        RECT 730.730 736.090 731.910 737.270 ;
        RECT 729.130 734.490 730.310 735.670 ;
        RECT 730.730 734.490 731.910 735.670 ;
        RECT 729.130 556.090 730.310 557.270 ;
        RECT 730.730 556.090 731.910 557.270 ;
        RECT 729.130 554.490 730.310 555.670 ;
        RECT 730.730 554.490 731.910 555.670 ;
        RECT 369.130 376.090 370.310 377.270 ;
        RECT 370.730 376.090 371.910 377.270 ;
        RECT 369.130 374.490 370.310 375.670 ;
        RECT 370.730 374.490 371.910 375.670 ;
        RECT 369.130 196.090 370.310 197.270 ;
        RECT 370.730 196.090 371.910 197.270 ;
        RECT 369.130 194.490 370.310 195.670 ;
        RECT 370.730 194.490 371.910 195.670 ;
        RECT 369.130 16.090 370.310 17.270 ;
        RECT 370.730 16.090 371.910 17.270 ;
        RECT 369.130 14.490 370.310 15.670 ;
        RECT 370.730 14.490 371.910 15.670 ;
        RECT 369.130 -2.910 370.310 -1.730 ;
        RECT 370.730 -2.910 371.910 -1.730 ;
        RECT 369.130 -4.510 370.310 -3.330 ;
        RECT 370.730 -4.510 371.910 -3.330 ;
        RECT 549.130 376.090 550.310 377.270 ;
        RECT 550.730 376.090 551.910 377.270 ;
        RECT 549.130 374.490 550.310 375.670 ;
        RECT 550.730 374.490 551.910 375.670 ;
        RECT 549.130 196.090 550.310 197.270 ;
        RECT 550.730 196.090 551.910 197.270 ;
        RECT 549.130 194.490 550.310 195.670 ;
        RECT 550.730 194.490 551.910 195.670 ;
        RECT 549.130 16.090 550.310 17.270 ;
        RECT 550.730 16.090 551.910 17.270 ;
        RECT 549.130 14.490 550.310 15.670 ;
        RECT 550.730 14.490 551.910 15.670 ;
        RECT 549.130 -2.910 550.310 -1.730 ;
        RECT 550.730 -2.910 551.910 -1.730 ;
        RECT 549.130 -4.510 550.310 -3.330 ;
        RECT 550.730 -4.510 551.910 -3.330 ;
        RECT 729.130 376.090 730.310 377.270 ;
        RECT 730.730 376.090 731.910 377.270 ;
        RECT 729.130 374.490 730.310 375.670 ;
        RECT 730.730 374.490 731.910 375.670 ;
        RECT 729.130 196.090 730.310 197.270 ;
        RECT 730.730 196.090 731.910 197.270 ;
        RECT 729.130 194.490 730.310 195.670 ;
        RECT 730.730 194.490 731.910 195.670 ;
        RECT 729.130 16.090 730.310 17.270 ;
        RECT 730.730 16.090 731.910 17.270 ;
        RECT 729.130 14.490 730.310 15.670 ;
        RECT 730.730 14.490 731.910 15.670 ;
        RECT 729.130 -2.910 730.310 -1.730 ;
        RECT 730.730 -2.910 731.910 -1.730 ;
        RECT 729.130 -4.510 730.310 -3.330 ;
        RECT 730.730 -4.510 731.910 -3.330 ;
        RECT 909.130 3523.010 910.310 3524.190 ;
        RECT 910.730 3523.010 911.910 3524.190 ;
        RECT 909.130 3521.410 910.310 3522.590 ;
        RECT 910.730 3521.410 911.910 3522.590 ;
        RECT 909.130 3436.090 910.310 3437.270 ;
        RECT 910.730 3436.090 911.910 3437.270 ;
        RECT 909.130 3434.490 910.310 3435.670 ;
        RECT 910.730 3434.490 911.910 3435.670 ;
        RECT 909.130 3256.090 910.310 3257.270 ;
        RECT 910.730 3256.090 911.910 3257.270 ;
        RECT 909.130 3254.490 910.310 3255.670 ;
        RECT 910.730 3254.490 911.910 3255.670 ;
        RECT 909.130 3076.090 910.310 3077.270 ;
        RECT 910.730 3076.090 911.910 3077.270 ;
        RECT 909.130 3074.490 910.310 3075.670 ;
        RECT 910.730 3074.490 911.910 3075.670 ;
        RECT 909.130 2896.090 910.310 2897.270 ;
        RECT 910.730 2896.090 911.910 2897.270 ;
        RECT 909.130 2894.490 910.310 2895.670 ;
        RECT 910.730 2894.490 911.910 2895.670 ;
        RECT 909.130 2716.090 910.310 2717.270 ;
        RECT 910.730 2716.090 911.910 2717.270 ;
        RECT 909.130 2714.490 910.310 2715.670 ;
        RECT 910.730 2714.490 911.910 2715.670 ;
        RECT 909.130 2536.090 910.310 2537.270 ;
        RECT 910.730 2536.090 911.910 2537.270 ;
        RECT 909.130 2534.490 910.310 2535.670 ;
        RECT 910.730 2534.490 911.910 2535.670 ;
        RECT 909.130 2356.090 910.310 2357.270 ;
        RECT 910.730 2356.090 911.910 2357.270 ;
        RECT 909.130 2354.490 910.310 2355.670 ;
        RECT 910.730 2354.490 911.910 2355.670 ;
        RECT 909.130 2176.090 910.310 2177.270 ;
        RECT 910.730 2176.090 911.910 2177.270 ;
        RECT 909.130 2174.490 910.310 2175.670 ;
        RECT 910.730 2174.490 911.910 2175.670 ;
        RECT 909.130 1996.090 910.310 1997.270 ;
        RECT 910.730 1996.090 911.910 1997.270 ;
        RECT 909.130 1994.490 910.310 1995.670 ;
        RECT 910.730 1994.490 911.910 1995.670 ;
        RECT 909.130 1816.090 910.310 1817.270 ;
        RECT 910.730 1816.090 911.910 1817.270 ;
        RECT 909.130 1814.490 910.310 1815.670 ;
        RECT 910.730 1814.490 911.910 1815.670 ;
        RECT 909.130 1636.090 910.310 1637.270 ;
        RECT 910.730 1636.090 911.910 1637.270 ;
        RECT 909.130 1634.490 910.310 1635.670 ;
        RECT 910.730 1634.490 911.910 1635.670 ;
        RECT 909.130 1456.090 910.310 1457.270 ;
        RECT 910.730 1456.090 911.910 1457.270 ;
        RECT 909.130 1454.490 910.310 1455.670 ;
        RECT 910.730 1454.490 911.910 1455.670 ;
        RECT 909.130 1276.090 910.310 1277.270 ;
        RECT 910.730 1276.090 911.910 1277.270 ;
        RECT 909.130 1274.490 910.310 1275.670 ;
        RECT 910.730 1274.490 911.910 1275.670 ;
        RECT 909.130 1096.090 910.310 1097.270 ;
        RECT 910.730 1096.090 911.910 1097.270 ;
        RECT 909.130 1094.490 910.310 1095.670 ;
        RECT 910.730 1094.490 911.910 1095.670 ;
        RECT 909.130 916.090 910.310 917.270 ;
        RECT 910.730 916.090 911.910 917.270 ;
        RECT 909.130 914.490 910.310 915.670 ;
        RECT 910.730 914.490 911.910 915.670 ;
        RECT 909.130 736.090 910.310 737.270 ;
        RECT 910.730 736.090 911.910 737.270 ;
        RECT 909.130 734.490 910.310 735.670 ;
        RECT 910.730 734.490 911.910 735.670 ;
        RECT 909.130 556.090 910.310 557.270 ;
        RECT 910.730 556.090 911.910 557.270 ;
        RECT 909.130 554.490 910.310 555.670 ;
        RECT 910.730 554.490 911.910 555.670 ;
        RECT 909.130 376.090 910.310 377.270 ;
        RECT 910.730 376.090 911.910 377.270 ;
        RECT 909.130 374.490 910.310 375.670 ;
        RECT 910.730 374.490 911.910 375.670 ;
        RECT 909.130 196.090 910.310 197.270 ;
        RECT 910.730 196.090 911.910 197.270 ;
        RECT 909.130 194.490 910.310 195.670 ;
        RECT 910.730 194.490 911.910 195.670 ;
        RECT 909.130 16.090 910.310 17.270 ;
        RECT 910.730 16.090 911.910 17.270 ;
        RECT 909.130 14.490 910.310 15.670 ;
        RECT 910.730 14.490 911.910 15.670 ;
        RECT 909.130 -2.910 910.310 -1.730 ;
        RECT 910.730 -2.910 911.910 -1.730 ;
        RECT 909.130 -4.510 910.310 -3.330 ;
        RECT 910.730 -4.510 911.910 -3.330 ;
        RECT 1089.130 3523.010 1090.310 3524.190 ;
        RECT 1090.730 3523.010 1091.910 3524.190 ;
        RECT 1089.130 3521.410 1090.310 3522.590 ;
        RECT 1090.730 3521.410 1091.910 3522.590 ;
        RECT 1089.130 3436.090 1090.310 3437.270 ;
        RECT 1090.730 3436.090 1091.910 3437.270 ;
        RECT 1089.130 3434.490 1090.310 3435.670 ;
        RECT 1090.730 3434.490 1091.910 3435.670 ;
        RECT 1089.130 3256.090 1090.310 3257.270 ;
        RECT 1090.730 3256.090 1091.910 3257.270 ;
        RECT 1089.130 3254.490 1090.310 3255.670 ;
        RECT 1090.730 3254.490 1091.910 3255.670 ;
        RECT 1089.130 3076.090 1090.310 3077.270 ;
        RECT 1090.730 3076.090 1091.910 3077.270 ;
        RECT 1089.130 3074.490 1090.310 3075.670 ;
        RECT 1090.730 3074.490 1091.910 3075.670 ;
        RECT 1089.130 2896.090 1090.310 2897.270 ;
        RECT 1090.730 2896.090 1091.910 2897.270 ;
        RECT 1089.130 2894.490 1090.310 2895.670 ;
        RECT 1090.730 2894.490 1091.910 2895.670 ;
        RECT 1089.130 2716.090 1090.310 2717.270 ;
        RECT 1090.730 2716.090 1091.910 2717.270 ;
        RECT 1089.130 2714.490 1090.310 2715.670 ;
        RECT 1090.730 2714.490 1091.910 2715.670 ;
        RECT 1089.130 2536.090 1090.310 2537.270 ;
        RECT 1090.730 2536.090 1091.910 2537.270 ;
        RECT 1089.130 2534.490 1090.310 2535.670 ;
        RECT 1090.730 2534.490 1091.910 2535.670 ;
        RECT 1089.130 2356.090 1090.310 2357.270 ;
        RECT 1090.730 2356.090 1091.910 2357.270 ;
        RECT 1089.130 2354.490 1090.310 2355.670 ;
        RECT 1090.730 2354.490 1091.910 2355.670 ;
        RECT 1089.130 2176.090 1090.310 2177.270 ;
        RECT 1090.730 2176.090 1091.910 2177.270 ;
        RECT 1089.130 2174.490 1090.310 2175.670 ;
        RECT 1090.730 2174.490 1091.910 2175.670 ;
        RECT 1089.130 1996.090 1090.310 1997.270 ;
        RECT 1090.730 1996.090 1091.910 1997.270 ;
        RECT 1089.130 1994.490 1090.310 1995.670 ;
        RECT 1090.730 1994.490 1091.910 1995.670 ;
        RECT 1089.130 1816.090 1090.310 1817.270 ;
        RECT 1090.730 1816.090 1091.910 1817.270 ;
        RECT 1089.130 1814.490 1090.310 1815.670 ;
        RECT 1090.730 1814.490 1091.910 1815.670 ;
        RECT 1089.130 1636.090 1090.310 1637.270 ;
        RECT 1090.730 1636.090 1091.910 1637.270 ;
        RECT 1089.130 1634.490 1090.310 1635.670 ;
        RECT 1090.730 1634.490 1091.910 1635.670 ;
        RECT 1089.130 1456.090 1090.310 1457.270 ;
        RECT 1090.730 1456.090 1091.910 1457.270 ;
        RECT 1089.130 1454.490 1090.310 1455.670 ;
        RECT 1090.730 1454.490 1091.910 1455.670 ;
        RECT 1089.130 1276.090 1090.310 1277.270 ;
        RECT 1090.730 1276.090 1091.910 1277.270 ;
        RECT 1089.130 1274.490 1090.310 1275.670 ;
        RECT 1090.730 1274.490 1091.910 1275.670 ;
        RECT 1089.130 1096.090 1090.310 1097.270 ;
        RECT 1090.730 1096.090 1091.910 1097.270 ;
        RECT 1089.130 1094.490 1090.310 1095.670 ;
        RECT 1090.730 1094.490 1091.910 1095.670 ;
        RECT 1089.130 916.090 1090.310 917.270 ;
        RECT 1090.730 916.090 1091.910 917.270 ;
        RECT 1089.130 914.490 1090.310 915.670 ;
        RECT 1090.730 914.490 1091.910 915.670 ;
        RECT 1089.130 736.090 1090.310 737.270 ;
        RECT 1090.730 736.090 1091.910 737.270 ;
        RECT 1089.130 734.490 1090.310 735.670 ;
        RECT 1090.730 734.490 1091.910 735.670 ;
        RECT 1089.130 556.090 1090.310 557.270 ;
        RECT 1090.730 556.090 1091.910 557.270 ;
        RECT 1089.130 554.490 1090.310 555.670 ;
        RECT 1090.730 554.490 1091.910 555.670 ;
        RECT 1089.130 376.090 1090.310 377.270 ;
        RECT 1090.730 376.090 1091.910 377.270 ;
        RECT 1089.130 374.490 1090.310 375.670 ;
        RECT 1090.730 374.490 1091.910 375.670 ;
        RECT 1089.130 196.090 1090.310 197.270 ;
        RECT 1090.730 196.090 1091.910 197.270 ;
        RECT 1089.130 194.490 1090.310 195.670 ;
        RECT 1090.730 194.490 1091.910 195.670 ;
        RECT 1089.130 16.090 1090.310 17.270 ;
        RECT 1090.730 16.090 1091.910 17.270 ;
        RECT 1089.130 14.490 1090.310 15.670 ;
        RECT 1090.730 14.490 1091.910 15.670 ;
        RECT 1089.130 -2.910 1090.310 -1.730 ;
        RECT 1090.730 -2.910 1091.910 -1.730 ;
        RECT 1089.130 -4.510 1090.310 -3.330 ;
        RECT 1090.730 -4.510 1091.910 -3.330 ;
        RECT 1269.130 3523.010 1270.310 3524.190 ;
        RECT 1270.730 3523.010 1271.910 3524.190 ;
        RECT 1269.130 3521.410 1270.310 3522.590 ;
        RECT 1270.730 3521.410 1271.910 3522.590 ;
        RECT 1269.130 3436.090 1270.310 3437.270 ;
        RECT 1270.730 3436.090 1271.910 3437.270 ;
        RECT 1269.130 3434.490 1270.310 3435.670 ;
        RECT 1270.730 3434.490 1271.910 3435.670 ;
        RECT 1269.130 3256.090 1270.310 3257.270 ;
        RECT 1270.730 3256.090 1271.910 3257.270 ;
        RECT 1269.130 3254.490 1270.310 3255.670 ;
        RECT 1270.730 3254.490 1271.910 3255.670 ;
        RECT 1269.130 3076.090 1270.310 3077.270 ;
        RECT 1270.730 3076.090 1271.910 3077.270 ;
        RECT 1269.130 3074.490 1270.310 3075.670 ;
        RECT 1270.730 3074.490 1271.910 3075.670 ;
        RECT 1269.130 2896.090 1270.310 2897.270 ;
        RECT 1270.730 2896.090 1271.910 2897.270 ;
        RECT 1269.130 2894.490 1270.310 2895.670 ;
        RECT 1270.730 2894.490 1271.910 2895.670 ;
        RECT 1269.130 2716.090 1270.310 2717.270 ;
        RECT 1270.730 2716.090 1271.910 2717.270 ;
        RECT 1269.130 2714.490 1270.310 2715.670 ;
        RECT 1270.730 2714.490 1271.910 2715.670 ;
        RECT 1269.130 2536.090 1270.310 2537.270 ;
        RECT 1270.730 2536.090 1271.910 2537.270 ;
        RECT 1269.130 2534.490 1270.310 2535.670 ;
        RECT 1270.730 2534.490 1271.910 2535.670 ;
        RECT 1269.130 2356.090 1270.310 2357.270 ;
        RECT 1270.730 2356.090 1271.910 2357.270 ;
        RECT 1269.130 2354.490 1270.310 2355.670 ;
        RECT 1270.730 2354.490 1271.910 2355.670 ;
        RECT 1269.130 2176.090 1270.310 2177.270 ;
        RECT 1270.730 2176.090 1271.910 2177.270 ;
        RECT 1269.130 2174.490 1270.310 2175.670 ;
        RECT 1270.730 2174.490 1271.910 2175.670 ;
        RECT 1269.130 1996.090 1270.310 1997.270 ;
        RECT 1270.730 1996.090 1271.910 1997.270 ;
        RECT 1269.130 1994.490 1270.310 1995.670 ;
        RECT 1270.730 1994.490 1271.910 1995.670 ;
        RECT 1269.130 1816.090 1270.310 1817.270 ;
        RECT 1270.730 1816.090 1271.910 1817.270 ;
        RECT 1269.130 1814.490 1270.310 1815.670 ;
        RECT 1270.730 1814.490 1271.910 1815.670 ;
        RECT 1269.130 1636.090 1270.310 1637.270 ;
        RECT 1270.730 1636.090 1271.910 1637.270 ;
        RECT 1269.130 1634.490 1270.310 1635.670 ;
        RECT 1270.730 1634.490 1271.910 1635.670 ;
        RECT 1269.130 1456.090 1270.310 1457.270 ;
        RECT 1270.730 1456.090 1271.910 1457.270 ;
        RECT 1269.130 1454.490 1270.310 1455.670 ;
        RECT 1270.730 1454.490 1271.910 1455.670 ;
        RECT 1269.130 1276.090 1270.310 1277.270 ;
        RECT 1270.730 1276.090 1271.910 1277.270 ;
        RECT 1269.130 1274.490 1270.310 1275.670 ;
        RECT 1270.730 1274.490 1271.910 1275.670 ;
        RECT 1269.130 1096.090 1270.310 1097.270 ;
        RECT 1270.730 1096.090 1271.910 1097.270 ;
        RECT 1269.130 1094.490 1270.310 1095.670 ;
        RECT 1270.730 1094.490 1271.910 1095.670 ;
        RECT 1269.130 916.090 1270.310 917.270 ;
        RECT 1270.730 916.090 1271.910 917.270 ;
        RECT 1269.130 914.490 1270.310 915.670 ;
        RECT 1270.730 914.490 1271.910 915.670 ;
        RECT 1269.130 736.090 1270.310 737.270 ;
        RECT 1270.730 736.090 1271.910 737.270 ;
        RECT 1269.130 734.490 1270.310 735.670 ;
        RECT 1270.730 734.490 1271.910 735.670 ;
        RECT 1269.130 556.090 1270.310 557.270 ;
        RECT 1270.730 556.090 1271.910 557.270 ;
        RECT 1269.130 554.490 1270.310 555.670 ;
        RECT 1270.730 554.490 1271.910 555.670 ;
        RECT 1269.130 376.090 1270.310 377.270 ;
        RECT 1270.730 376.090 1271.910 377.270 ;
        RECT 1269.130 374.490 1270.310 375.670 ;
        RECT 1270.730 374.490 1271.910 375.670 ;
        RECT 1269.130 196.090 1270.310 197.270 ;
        RECT 1270.730 196.090 1271.910 197.270 ;
        RECT 1269.130 194.490 1270.310 195.670 ;
        RECT 1270.730 194.490 1271.910 195.670 ;
        RECT 1269.130 16.090 1270.310 17.270 ;
        RECT 1270.730 16.090 1271.910 17.270 ;
        RECT 1269.130 14.490 1270.310 15.670 ;
        RECT 1270.730 14.490 1271.910 15.670 ;
        RECT 1269.130 -2.910 1270.310 -1.730 ;
        RECT 1270.730 -2.910 1271.910 -1.730 ;
        RECT 1269.130 -4.510 1270.310 -3.330 ;
        RECT 1270.730 -4.510 1271.910 -3.330 ;
        RECT 1449.130 3523.010 1450.310 3524.190 ;
        RECT 1450.730 3523.010 1451.910 3524.190 ;
        RECT 1449.130 3521.410 1450.310 3522.590 ;
        RECT 1450.730 3521.410 1451.910 3522.590 ;
        RECT 1449.130 3436.090 1450.310 3437.270 ;
        RECT 1450.730 3436.090 1451.910 3437.270 ;
        RECT 1449.130 3434.490 1450.310 3435.670 ;
        RECT 1450.730 3434.490 1451.910 3435.670 ;
        RECT 1449.130 3256.090 1450.310 3257.270 ;
        RECT 1450.730 3256.090 1451.910 3257.270 ;
        RECT 1449.130 3254.490 1450.310 3255.670 ;
        RECT 1450.730 3254.490 1451.910 3255.670 ;
        RECT 1449.130 3076.090 1450.310 3077.270 ;
        RECT 1450.730 3076.090 1451.910 3077.270 ;
        RECT 1449.130 3074.490 1450.310 3075.670 ;
        RECT 1450.730 3074.490 1451.910 3075.670 ;
        RECT 1449.130 2896.090 1450.310 2897.270 ;
        RECT 1450.730 2896.090 1451.910 2897.270 ;
        RECT 1449.130 2894.490 1450.310 2895.670 ;
        RECT 1450.730 2894.490 1451.910 2895.670 ;
        RECT 1449.130 2716.090 1450.310 2717.270 ;
        RECT 1450.730 2716.090 1451.910 2717.270 ;
        RECT 1449.130 2714.490 1450.310 2715.670 ;
        RECT 1450.730 2714.490 1451.910 2715.670 ;
        RECT 1449.130 2536.090 1450.310 2537.270 ;
        RECT 1450.730 2536.090 1451.910 2537.270 ;
        RECT 1449.130 2534.490 1450.310 2535.670 ;
        RECT 1450.730 2534.490 1451.910 2535.670 ;
        RECT 1449.130 2356.090 1450.310 2357.270 ;
        RECT 1450.730 2356.090 1451.910 2357.270 ;
        RECT 1449.130 2354.490 1450.310 2355.670 ;
        RECT 1450.730 2354.490 1451.910 2355.670 ;
        RECT 1449.130 2176.090 1450.310 2177.270 ;
        RECT 1450.730 2176.090 1451.910 2177.270 ;
        RECT 1449.130 2174.490 1450.310 2175.670 ;
        RECT 1450.730 2174.490 1451.910 2175.670 ;
        RECT 1449.130 1996.090 1450.310 1997.270 ;
        RECT 1450.730 1996.090 1451.910 1997.270 ;
        RECT 1449.130 1994.490 1450.310 1995.670 ;
        RECT 1450.730 1994.490 1451.910 1995.670 ;
        RECT 1449.130 1816.090 1450.310 1817.270 ;
        RECT 1450.730 1816.090 1451.910 1817.270 ;
        RECT 1449.130 1814.490 1450.310 1815.670 ;
        RECT 1450.730 1814.490 1451.910 1815.670 ;
        RECT 1449.130 1636.090 1450.310 1637.270 ;
        RECT 1450.730 1636.090 1451.910 1637.270 ;
        RECT 1449.130 1634.490 1450.310 1635.670 ;
        RECT 1450.730 1634.490 1451.910 1635.670 ;
        RECT 1449.130 1456.090 1450.310 1457.270 ;
        RECT 1450.730 1456.090 1451.910 1457.270 ;
        RECT 1449.130 1454.490 1450.310 1455.670 ;
        RECT 1450.730 1454.490 1451.910 1455.670 ;
        RECT 1449.130 1276.090 1450.310 1277.270 ;
        RECT 1450.730 1276.090 1451.910 1277.270 ;
        RECT 1449.130 1274.490 1450.310 1275.670 ;
        RECT 1450.730 1274.490 1451.910 1275.670 ;
        RECT 1449.130 1096.090 1450.310 1097.270 ;
        RECT 1450.730 1096.090 1451.910 1097.270 ;
        RECT 1449.130 1094.490 1450.310 1095.670 ;
        RECT 1450.730 1094.490 1451.910 1095.670 ;
        RECT 1449.130 916.090 1450.310 917.270 ;
        RECT 1450.730 916.090 1451.910 917.270 ;
        RECT 1449.130 914.490 1450.310 915.670 ;
        RECT 1450.730 914.490 1451.910 915.670 ;
        RECT 1449.130 736.090 1450.310 737.270 ;
        RECT 1450.730 736.090 1451.910 737.270 ;
        RECT 1449.130 734.490 1450.310 735.670 ;
        RECT 1450.730 734.490 1451.910 735.670 ;
        RECT 1449.130 556.090 1450.310 557.270 ;
        RECT 1450.730 556.090 1451.910 557.270 ;
        RECT 1449.130 554.490 1450.310 555.670 ;
        RECT 1450.730 554.490 1451.910 555.670 ;
        RECT 1449.130 376.090 1450.310 377.270 ;
        RECT 1450.730 376.090 1451.910 377.270 ;
        RECT 1449.130 374.490 1450.310 375.670 ;
        RECT 1450.730 374.490 1451.910 375.670 ;
        RECT 1449.130 196.090 1450.310 197.270 ;
        RECT 1450.730 196.090 1451.910 197.270 ;
        RECT 1449.130 194.490 1450.310 195.670 ;
        RECT 1450.730 194.490 1451.910 195.670 ;
        RECT 1449.130 16.090 1450.310 17.270 ;
        RECT 1450.730 16.090 1451.910 17.270 ;
        RECT 1449.130 14.490 1450.310 15.670 ;
        RECT 1450.730 14.490 1451.910 15.670 ;
        RECT 1449.130 -2.910 1450.310 -1.730 ;
        RECT 1450.730 -2.910 1451.910 -1.730 ;
        RECT 1449.130 -4.510 1450.310 -3.330 ;
        RECT 1450.730 -4.510 1451.910 -3.330 ;
        RECT 1629.130 3523.010 1630.310 3524.190 ;
        RECT 1630.730 3523.010 1631.910 3524.190 ;
        RECT 1629.130 3521.410 1630.310 3522.590 ;
        RECT 1630.730 3521.410 1631.910 3522.590 ;
        RECT 1629.130 3436.090 1630.310 3437.270 ;
        RECT 1630.730 3436.090 1631.910 3437.270 ;
        RECT 1629.130 3434.490 1630.310 3435.670 ;
        RECT 1630.730 3434.490 1631.910 3435.670 ;
        RECT 1629.130 3256.090 1630.310 3257.270 ;
        RECT 1630.730 3256.090 1631.910 3257.270 ;
        RECT 1629.130 3254.490 1630.310 3255.670 ;
        RECT 1630.730 3254.490 1631.910 3255.670 ;
        RECT 1629.130 3076.090 1630.310 3077.270 ;
        RECT 1630.730 3076.090 1631.910 3077.270 ;
        RECT 1629.130 3074.490 1630.310 3075.670 ;
        RECT 1630.730 3074.490 1631.910 3075.670 ;
        RECT 1629.130 2896.090 1630.310 2897.270 ;
        RECT 1630.730 2896.090 1631.910 2897.270 ;
        RECT 1629.130 2894.490 1630.310 2895.670 ;
        RECT 1630.730 2894.490 1631.910 2895.670 ;
        RECT 1629.130 2716.090 1630.310 2717.270 ;
        RECT 1630.730 2716.090 1631.910 2717.270 ;
        RECT 1629.130 2714.490 1630.310 2715.670 ;
        RECT 1630.730 2714.490 1631.910 2715.670 ;
        RECT 1629.130 2536.090 1630.310 2537.270 ;
        RECT 1630.730 2536.090 1631.910 2537.270 ;
        RECT 1629.130 2534.490 1630.310 2535.670 ;
        RECT 1630.730 2534.490 1631.910 2535.670 ;
        RECT 1629.130 2356.090 1630.310 2357.270 ;
        RECT 1630.730 2356.090 1631.910 2357.270 ;
        RECT 1629.130 2354.490 1630.310 2355.670 ;
        RECT 1630.730 2354.490 1631.910 2355.670 ;
        RECT 1629.130 2176.090 1630.310 2177.270 ;
        RECT 1630.730 2176.090 1631.910 2177.270 ;
        RECT 1629.130 2174.490 1630.310 2175.670 ;
        RECT 1630.730 2174.490 1631.910 2175.670 ;
        RECT 1629.130 1996.090 1630.310 1997.270 ;
        RECT 1630.730 1996.090 1631.910 1997.270 ;
        RECT 1629.130 1994.490 1630.310 1995.670 ;
        RECT 1630.730 1994.490 1631.910 1995.670 ;
        RECT 1629.130 1816.090 1630.310 1817.270 ;
        RECT 1630.730 1816.090 1631.910 1817.270 ;
        RECT 1629.130 1814.490 1630.310 1815.670 ;
        RECT 1630.730 1814.490 1631.910 1815.670 ;
        RECT 1629.130 1636.090 1630.310 1637.270 ;
        RECT 1630.730 1636.090 1631.910 1637.270 ;
        RECT 1629.130 1634.490 1630.310 1635.670 ;
        RECT 1630.730 1634.490 1631.910 1635.670 ;
        RECT 1629.130 1456.090 1630.310 1457.270 ;
        RECT 1630.730 1456.090 1631.910 1457.270 ;
        RECT 1629.130 1454.490 1630.310 1455.670 ;
        RECT 1630.730 1454.490 1631.910 1455.670 ;
        RECT 1629.130 1276.090 1630.310 1277.270 ;
        RECT 1630.730 1276.090 1631.910 1277.270 ;
        RECT 1629.130 1274.490 1630.310 1275.670 ;
        RECT 1630.730 1274.490 1631.910 1275.670 ;
        RECT 1629.130 1096.090 1630.310 1097.270 ;
        RECT 1630.730 1096.090 1631.910 1097.270 ;
        RECT 1629.130 1094.490 1630.310 1095.670 ;
        RECT 1630.730 1094.490 1631.910 1095.670 ;
        RECT 1629.130 916.090 1630.310 917.270 ;
        RECT 1630.730 916.090 1631.910 917.270 ;
        RECT 1629.130 914.490 1630.310 915.670 ;
        RECT 1630.730 914.490 1631.910 915.670 ;
        RECT 1629.130 736.090 1630.310 737.270 ;
        RECT 1630.730 736.090 1631.910 737.270 ;
        RECT 1629.130 734.490 1630.310 735.670 ;
        RECT 1630.730 734.490 1631.910 735.670 ;
        RECT 1629.130 556.090 1630.310 557.270 ;
        RECT 1630.730 556.090 1631.910 557.270 ;
        RECT 1629.130 554.490 1630.310 555.670 ;
        RECT 1630.730 554.490 1631.910 555.670 ;
        RECT 1629.130 376.090 1630.310 377.270 ;
        RECT 1630.730 376.090 1631.910 377.270 ;
        RECT 1629.130 374.490 1630.310 375.670 ;
        RECT 1630.730 374.490 1631.910 375.670 ;
        RECT 1629.130 196.090 1630.310 197.270 ;
        RECT 1630.730 196.090 1631.910 197.270 ;
        RECT 1629.130 194.490 1630.310 195.670 ;
        RECT 1630.730 194.490 1631.910 195.670 ;
        RECT 1629.130 16.090 1630.310 17.270 ;
        RECT 1630.730 16.090 1631.910 17.270 ;
        RECT 1629.130 14.490 1630.310 15.670 ;
        RECT 1630.730 14.490 1631.910 15.670 ;
        RECT 1629.130 -2.910 1630.310 -1.730 ;
        RECT 1630.730 -2.910 1631.910 -1.730 ;
        RECT 1629.130 -4.510 1630.310 -3.330 ;
        RECT 1630.730 -4.510 1631.910 -3.330 ;
        RECT 1809.130 3523.010 1810.310 3524.190 ;
        RECT 1810.730 3523.010 1811.910 3524.190 ;
        RECT 1809.130 3521.410 1810.310 3522.590 ;
        RECT 1810.730 3521.410 1811.910 3522.590 ;
        RECT 1809.130 3436.090 1810.310 3437.270 ;
        RECT 1810.730 3436.090 1811.910 3437.270 ;
        RECT 1809.130 3434.490 1810.310 3435.670 ;
        RECT 1810.730 3434.490 1811.910 3435.670 ;
        RECT 1809.130 3256.090 1810.310 3257.270 ;
        RECT 1810.730 3256.090 1811.910 3257.270 ;
        RECT 1809.130 3254.490 1810.310 3255.670 ;
        RECT 1810.730 3254.490 1811.910 3255.670 ;
        RECT 1809.130 3076.090 1810.310 3077.270 ;
        RECT 1810.730 3076.090 1811.910 3077.270 ;
        RECT 1809.130 3074.490 1810.310 3075.670 ;
        RECT 1810.730 3074.490 1811.910 3075.670 ;
        RECT 1809.130 2896.090 1810.310 2897.270 ;
        RECT 1810.730 2896.090 1811.910 2897.270 ;
        RECT 1809.130 2894.490 1810.310 2895.670 ;
        RECT 1810.730 2894.490 1811.910 2895.670 ;
        RECT 1809.130 2716.090 1810.310 2717.270 ;
        RECT 1810.730 2716.090 1811.910 2717.270 ;
        RECT 1809.130 2714.490 1810.310 2715.670 ;
        RECT 1810.730 2714.490 1811.910 2715.670 ;
        RECT 1809.130 2536.090 1810.310 2537.270 ;
        RECT 1810.730 2536.090 1811.910 2537.270 ;
        RECT 1809.130 2534.490 1810.310 2535.670 ;
        RECT 1810.730 2534.490 1811.910 2535.670 ;
        RECT 1809.130 2356.090 1810.310 2357.270 ;
        RECT 1810.730 2356.090 1811.910 2357.270 ;
        RECT 1809.130 2354.490 1810.310 2355.670 ;
        RECT 1810.730 2354.490 1811.910 2355.670 ;
        RECT 1809.130 2176.090 1810.310 2177.270 ;
        RECT 1810.730 2176.090 1811.910 2177.270 ;
        RECT 1809.130 2174.490 1810.310 2175.670 ;
        RECT 1810.730 2174.490 1811.910 2175.670 ;
        RECT 1809.130 1996.090 1810.310 1997.270 ;
        RECT 1810.730 1996.090 1811.910 1997.270 ;
        RECT 1809.130 1994.490 1810.310 1995.670 ;
        RECT 1810.730 1994.490 1811.910 1995.670 ;
        RECT 1809.130 1816.090 1810.310 1817.270 ;
        RECT 1810.730 1816.090 1811.910 1817.270 ;
        RECT 1809.130 1814.490 1810.310 1815.670 ;
        RECT 1810.730 1814.490 1811.910 1815.670 ;
        RECT 1809.130 1636.090 1810.310 1637.270 ;
        RECT 1810.730 1636.090 1811.910 1637.270 ;
        RECT 1809.130 1634.490 1810.310 1635.670 ;
        RECT 1810.730 1634.490 1811.910 1635.670 ;
        RECT 1809.130 1456.090 1810.310 1457.270 ;
        RECT 1810.730 1456.090 1811.910 1457.270 ;
        RECT 1809.130 1454.490 1810.310 1455.670 ;
        RECT 1810.730 1454.490 1811.910 1455.670 ;
        RECT 1809.130 1276.090 1810.310 1277.270 ;
        RECT 1810.730 1276.090 1811.910 1277.270 ;
        RECT 1809.130 1274.490 1810.310 1275.670 ;
        RECT 1810.730 1274.490 1811.910 1275.670 ;
        RECT 1809.130 1096.090 1810.310 1097.270 ;
        RECT 1810.730 1096.090 1811.910 1097.270 ;
        RECT 1809.130 1094.490 1810.310 1095.670 ;
        RECT 1810.730 1094.490 1811.910 1095.670 ;
        RECT 1809.130 916.090 1810.310 917.270 ;
        RECT 1810.730 916.090 1811.910 917.270 ;
        RECT 1809.130 914.490 1810.310 915.670 ;
        RECT 1810.730 914.490 1811.910 915.670 ;
        RECT 1809.130 736.090 1810.310 737.270 ;
        RECT 1810.730 736.090 1811.910 737.270 ;
        RECT 1809.130 734.490 1810.310 735.670 ;
        RECT 1810.730 734.490 1811.910 735.670 ;
        RECT 1809.130 556.090 1810.310 557.270 ;
        RECT 1810.730 556.090 1811.910 557.270 ;
        RECT 1809.130 554.490 1810.310 555.670 ;
        RECT 1810.730 554.490 1811.910 555.670 ;
        RECT 1809.130 376.090 1810.310 377.270 ;
        RECT 1810.730 376.090 1811.910 377.270 ;
        RECT 1809.130 374.490 1810.310 375.670 ;
        RECT 1810.730 374.490 1811.910 375.670 ;
        RECT 1809.130 196.090 1810.310 197.270 ;
        RECT 1810.730 196.090 1811.910 197.270 ;
        RECT 1809.130 194.490 1810.310 195.670 ;
        RECT 1810.730 194.490 1811.910 195.670 ;
        RECT 1809.130 16.090 1810.310 17.270 ;
        RECT 1810.730 16.090 1811.910 17.270 ;
        RECT 1809.130 14.490 1810.310 15.670 ;
        RECT 1810.730 14.490 1811.910 15.670 ;
        RECT 1809.130 -2.910 1810.310 -1.730 ;
        RECT 1810.730 -2.910 1811.910 -1.730 ;
        RECT 1809.130 -4.510 1810.310 -3.330 ;
        RECT 1810.730 -4.510 1811.910 -3.330 ;
        RECT 1989.130 3523.010 1990.310 3524.190 ;
        RECT 1990.730 3523.010 1991.910 3524.190 ;
        RECT 1989.130 3521.410 1990.310 3522.590 ;
        RECT 1990.730 3521.410 1991.910 3522.590 ;
        RECT 1989.130 3436.090 1990.310 3437.270 ;
        RECT 1990.730 3436.090 1991.910 3437.270 ;
        RECT 1989.130 3434.490 1990.310 3435.670 ;
        RECT 1990.730 3434.490 1991.910 3435.670 ;
        RECT 1989.130 3256.090 1990.310 3257.270 ;
        RECT 1990.730 3256.090 1991.910 3257.270 ;
        RECT 1989.130 3254.490 1990.310 3255.670 ;
        RECT 1990.730 3254.490 1991.910 3255.670 ;
        RECT 1989.130 3076.090 1990.310 3077.270 ;
        RECT 1990.730 3076.090 1991.910 3077.270 ;
        RECT 1989.130 3074.490 1990.310 3075.670 ;
        RECT 1990.730 3074.490 1991.910 3075.670 ;
        RECT 1989.130 2896.090 1990.310 2897.270 ;
        RECT 1990.730 2896.090 1991.910 2897.270 ;
        RECT 1989.130 2894.490 1990.310 2895.670 ;
        RECT 1990.730 2894.490 1991.910 2895.670 ;
        RECT 1989.130 2716.090 1990.310 2717.270 ;
        RECT 1990.730 2716.090 1991.910 2717.270 ;
        RECT 1989.130 2714.490 1990.310 2715.670 ;
        RECT 1990.730 2714.490 1991.910 2715.670 ;
        RECT 1989.130 2536.090 1990.310 2537.270 ;
        RECT 1990.730 2536.090 1991.910 2537.270 ;
        RECT 1989.130 2534.490 1990.310 2535.670 ;
        RECT 1990.730 2534.490 1991.910 2535.670 ;
        RECT 1989.130 2356.090 1990.310 2357.270 ;
        RECT 1990.730 2356.090 1991.910 2357.270 ;
        RECT 1989.130 2354.490 1990.310 2355.670 ;
        RECT 1990.730 2354.490 1991.910 2355.670 ;
        RECT 1989.130 2176.090 1990.310 2177.270 ;
        RECT 1990.730 2176.090 1991.910 2177.270 ;
        RECT 1989.130 2174.490 1990.310 2175.670 ;
        RECT 1990.730 2174.490 1991.910 2175.670 ;
        RECT 1989.130 1996.090 1990.310 1997.270 ;
        RECT 1990.730 1996.090 1991.910 1997.270 ;
        RECT 1989.130 1994.490 1990.310 1995.670 ;
        RECT 1990.730 1994.490 1991.910 1995.670 ;
        RECT 1989.130 1816.090 1990.310 1817.270 ;
        RECT 1990.730 1816.090 1991.910 1817.270 ;
        RECT 1989.130 1814.490 1990.310 1815.670 ;
        RECT 1990.730 1814.490 1991.910 1815.670 ;
        RECT 1989.130 1636.090 1990.310 1637.270 ;
        RECT 1990.730 1636.090 1991.910 1637.270 ;
        RECT 1989.130 1634.490 1990.310 1635.670 ;
        RECT 1990.730 1634.490 1991.910 1635.670 ;
        RECT 1989.130 1456.090 1990.310 1457.270 ;
        RECT 1990.730 1456.090 1991.910 1457.270 ;
        RECT 1989.130 1454.490 1990.310 1455.670 ;
        RECT 1990.730 1454.490 1991.910 1455.670 ;
        RECT 1989.130 1276.090 1990.310 1277.270 ;
        RECT 1990.730 1276.090 1991.910 1277.270 ;
        RECT 1989.130 1274.490 1990.310 1275.670 ;
        RECT 1990.730 1274.490 1991.910 1275.670 ;
        RECT 1989.130 1096.090 1990.310 1097.270 ;
        RECT 1990.730 1096.090 1991.910 1097.270 ;
        RECT 1989.130 1094.490 1990.310 1095.670 ;
        RECT 1990.730 1094.490 1991.910 1095.670 ;
        RECT 1989.130 916.090 1990.310 917.270 ;
        RECT 1990.730 916.090 1991.910 917.270 ;
        RECT 1989.130 914.490 1990.310 915.670 ;
        RECT 1990.730 914.490 1991.910 915.670 ;
        RECT 1989.130 736.090 1990.310 737.270 ;
        RECT 1990.730 736.090 1991.910 737.270 ;
        RECT 1989.130 734.490 1990.310 735.670 ;
        RECT 1990.730 734.490 1991.910 735.670 ;
        RECT 1989.130 556.090 1990.310 557.270 ;
        RECT 1990.730 556.090 1991.910 557.270 ;
        RECT 1989.130 554.490 1990.310 555.670 ;
        RECT 1990.730 554.490 1991.910 555.670 ;
        RECT 1989.130 376.090 1990.310 377.270 ;
        RECT 1990.730 376.090 1991.910 377.270 ;
        RECT 1989.130 374.490 1990.310 375.670 ;
        RECT 1990.730 374.490 1991.910 375.670 ;
        RECT 1989.130 196.090 1990.310 197.270 ;
        RECT 1990.730 196.090 1991.910 197.270 ;
        RECT 1989.130 194.490 1990.310 195.670 ;
        RECT 1990.730 194.490 1991.910 195.670 ;
        RECT 1989.130 16.090 1990.310 17.270 ;
        RECT 1990.730 16.090 1991.910 17.270 ;
        RECT 1989.130 14.490 1990.310 15.670 ;
        RECT 1990.730 14.490 1991.910 15.670 ;
        RECT 1989.130 -2.910 1990.310 -1.730 ;
        RECT 1990.730 -2.910 1991.910 -1.730 ;
        RECT 1989.130 -4.510 1990.310 -3.330 ;
        RECT 1990.730 -4.510 1991.910 -3.330 ;
        RECT 2169.130 3523.010 2170.310 3524.190 ;
        RECT 2170.730 3523.010 2171.910 3524.190 ;
        RECT 2169.130 3521.410 2170.310 3522.590 ;
        RECT 2170.730 3521.410 2171.910 3522.590 ;
        RECT 2169.130 3436.090 2170.310 3437.270 ;
        RECT 2170.730 3436.090 2171.910 3437.270 ;
        RECT 2169.130 3434.490 2170.310 3435.670 ;
        RECT 2170.730 3434.490 2171.910 3435.670 ;
        RECT 2169.130 3256.090 2170.310 3257.270 ;
        RECT 2170.730 3256.090 2171.910 3257.270 ;
        RECT 2169.130 3254.490 2170.310 3255.670 ;
        RECT 2170.730 3254.490 2171.910 3255.670 ;
        RECT 2169.130 3076.090 2170.310 3077.270 ;
        RECT 2170.730 3076.090 2171.910 3077.270 ;
        RECT 2169.130 3074.490 2170.310 3075.670 ;
        RECT 2170.730 3074.490 2171.910 3075.670 ;
        RECT 2169.130 2896.090 2170.310 2897.270 ;
        RECT 2170.730 2896.090 2171.910 2897.270 ;
        RECT 2169.130 2894.490 2170.310 2895.670 ;
        RECT 2170.730 2894.490 2171.910 2895.670 ;
        RECT 2169.130 2716.090 2170.310 2717.270 ;
        RECT 2170.730 2716.090 2171.910 2717.270 ;
        RECT 2169.130 2714.490 2170.310 2715.670 ;
        RECT 2170.730 2714.490 2171.910 2715.670 ;
        RECT 2169.130 2536.090 2170.310 2537.270 ;
        RECT 2170.730 2536.090 2171.910 2537.270 ;
        RECT 2169.130 2534.490 2170.310 2535.670 ;
        RECT 2170.730 2534.490 2171.910 2535.670 ;
        RECT 2169.130 2356.090 2170.310 2357.270 ;
        RECT 2170.730 2356.090 2171.910 2357.270 ;
        RECT 2169.130 2354.490 2170.310 2355.670 ;
        RECT 2170.730 2354.490 2171.910 2355.670 ;
        RECT 2169.130 2176.090 2170.310 2177.270 ;
        RECT 2170.730 2176.090 2171.910 2177.270 ;
        RECT 2169.130 2174.490 2170.310 2175.670 ;
        RECT 2170.730 2174.490 2171.910 2175.670 ;
        RECT 2169.130 1996.090 2170.310 1997.270 ;
        RECT 2170.730 1996.090 2171.910 1997.270 ;
        RECT 2169.130 1994.490 2170.310 1995.670 ;
        RECT 2170.730 1994.490 2171.910 1995.670 ;
        RECT 2169.130 1816.090 2170.310 1817.270 ;
        RECT 2170.730 1816.090 2171.910 1817.270 ;
        RECT 2169.130 1814.490 2170.310 1815.670 ;
        RECT 2170.730 1814.490 2171.910 1815.670 ;
        RECT 2169.130 1636.090 2170.310 1637.270 ;
        RECT 2170.730 1636.090 2171.910 1637.270 ;
        RECT 2169.130 1634.490 2170.310 1635.670 ;
        RECT 2170.730 1634.490 2171.910 1635.670 ;
        RECT 2169.130 1456.090 2170.310 1457.270 ;
        RECT 2170.730 1456.090 2171.910 1457.270 ;
        RECT 2169.130 1454.490 2170.310 1455.670 ;
        RECT 2170.730 1454.490 2171.910 1455.670 ;
        RECT 2169.130 1276.090 2170.310 1277.270 ;
        RECT 2170.730 1276.090 2171.910 1277.270 ;
        RECT 2169.130 1274.490 2170.310 1275.670 ;
        RECT 2170.730 1274.490 2171.910 1275.670 ;
        RECT 2169.130 1096.090 2170.310 1097.270 ;
        RECT 2170.730 1096.090 2171.910 1097.270 ;
        RECT 2169.130 1094.490 2170.310 1095.670 ;
        RECT 2170.730 1094.490 2171.910 1095.670 ;
        RECT 2169.130 916.090 2170.310 917.270 ;
        RECT 2170.730 916.090 2171.910 917.270 ;
        RECT 2169.130 914.490 2170.310 915.670 ;
        RECT 2170.730 914.490 2171.910 915.670 ;
        RECT 2169.130 736.090 2170.310 737.270 ;
        RECT 2170.730 736.090 2171.910 737.270 ;
        RECT 2169.130 734.490 2170.310 735.670 ;
        RECT 2170.730 734.490 2171.910 735.670 ;
        RECT 2169.130 556.090 2170.310 557.270 ;
        RECT 2170.730 556.090 2171.910 557.270 ;
        RECT 2169.130 554.490 2170.310 555.670 ;
        RECT 2170.730 554.490 2171.910 555.670 ;
        RECT 2169.130 376.090 2170.310 377.270 ;
        RECT 2170.730 376.090 2171.910 377.270 ;
        RECT 2169.130 374.490 2170.310 375.670 ;
        RECT 2170.730 374.490 2171.910 375.670 ;
        RECT 2169.130 196.090 2170.310 197.270 ;
        RECT 2170.730 196.090 2171.910 197.270 ;
        RECT 2169.130 194.490 2170.310 195.670 ;
        RECT 2170.730 194.490 2171.910 195.670 ;
        RECT 2169.130 16.090 2170.310 17.270 ;
        RECT 2170.730 16.090 2171.910 17.270 ;
        RECT 2169.130 14.490 2170.310 15.670 ;
        RECT 2170.730 14.490 2171.910 15.670 ;
        RECT 2169.130 -2.910 2170.310 -1.730 ;
        RECT 2170.730 -2.910 2171.910 -1.730 ;
        RECT 2169.130 -4.510 2170.310 -3.330 ;
        RECT 2170.730 -4.510 2171.910 -3.330 ;
        RECT 2349.130 3523.010 2350.310 3524.190 ;
        RECT 2350.730 3523.010 2351.910 3524.190 ;
        RECT 2349.130 3521.410 2350.310 3522.590 ;
        RECT 2350.730 3521.410 2351.910 3522.590 ;
        RECT 2349.130 3436.090 2350.310 3437.270 ;
        RECT 2350.730 3436.090 2351.910 3437.270 ;
        RECT 2349.130 3434.490 2350.310 3435.670 ;
        RECT 2350.730 3434.490 2351.910 3435.670 ;
        RECT 2349.130 3256.090 2350.310 3257.270 ;
        RECT 2350.730 3256.090 2351.910 3257.270 ;
        RECT 2349.130 3254.490 2350.310 3255.670 ;
        RECT 2350.730 3254.490 2351.910 3255.670 ;
        RECT 2349.130 3076.090 2350.310 3077.270 ;
        RECT 2350.730 3076.090 2351.910 3077.270 ;
        RECT 2349.130 3074.490 2350.310 3075.670 ;
        RECT 2350.730 3074.490 2351.910 3075.670 ;
        RECT 2349.130 2896.090 2350.310 2897.270 ;
        RECT 2350.730 2896.090 2351.910 2897.270 ;
        RECT 2349.130 2894.490 2350.310 2895.670 ;
        RECT 2350.730 2894.490 2351.910 2895.670 ;
        RECT 2349.130 2716.090 2350.310 2717.270 ;
        RECT 2350.730 2716.090 2351.910 2717.270 ;
        RECT 2349.130 2714.490 2350.310 2715.670 ;
        RECT 2350.730 2714.490 2351.910 2715.670 ;
        RECT 2349.130 2536.090 2350.310 2537.270 ;
        RECT 2350.730 2536.090 2351.910 2537.270 ;
        RECT 2349.130 2534.490 2350.310 2535.670 ;
        RECT 2350.730 2534.490 2351.910 2535.670 ;
        RECT 2349.130 2356.090 2350.310 2357.270 ;
        RECT 2350.730 2356.090 2351.910 2357.270 ;
        RECT 2349.130 2354.490 2350.310 2355.670 ;
        RECT 2350.730 2354.490 2351.910 2355.670 ;
        RECT 2349.130 2176.090 2350.310 2177.270 ;
        RECT 2350.730 2176.090 2351.910 2177.270 ;
        RECT 2349.130 2174.490 2350.310 2175.670 ;
        RECT 2350.730 2174.490 2351.910 2175.670 ;
        RECT 2349.130 1996.090 2350.310 1997.270 ;
        RECT 2350.730 1996.090 2351.910 1997.270 ;
        RECT 2349.130 1994.490 2350.310 1995.670 ;
        RECT 2350.730 1994.490 2351.910 1995.670 ;
        RECT 2349.130 1816.090 2350.310 1817.270 ;
        RECT 2350.730 1816.090 2351.910 1817.270 ;
        RECT 2349.130 1814.490 2350.310 1815.670 ;
        RECT 2350.730 1814.490 2351.910 1815.670 ;
        RECT 2349.130 1636.090 2350.310 1637.270 ;
        RECT 2350.730 1636.090 2351.910 1637.270 ;
        RECT 2349.130 1634.490 2350.310 1635.670 ;
        RECT 2350.730 1634.490 2351.910 1635.670 ;
        RECT 2349.130 1456.090 2350.310 1457.270 ;
        RECT 2350.730 1456.090 2351.910 1457.270 ;
        RECT 2349.130 1454.490 2350.310 1455.670 ;
        RECT 2350.730 1454.490 2351.910 1455.670 ;
        RECT 2349.130 1276.090 2350.310 1277.270 ;
        RECT 2350.730 1276.090 2351.910 1277.270 ;
        RECT 2349.130 1274.490 2350.310 1275.670 ;
        RECT 2350.730 1274.490 2351.910 1275.670 ;
        RECT 2349.130 1096.090 2350.310 1097.270 ;
        RECT 2350.730 1096.090 2351.910 1097.270 ;
        RECT 2349.130 1094.490 2350.310 1095.670 ;
        RECT 2350.730 1094.490 2351.910 1095.670 ;
        RECT 2349.130 916.090 2350.310 917.270 ;
        RECT 2350.730 916.090 2351.910 917.270 ;
        RECT 2349.130 914.490 2350.310 915.670 ;
        RECT 2350.730 914.490 2351.910 915.670 ;
        RECT 2349.130 736.090 2350.310 737.270 ;
        RECT 2350.730 736.090 2351.910 737.270 ;
        RECT 2349.130 734.490 2350.310 735.670 ;
        RECT 2350.730 734.490 2351.910 735.670 ;
        RECT 2349.130 556.090 2350.310 557.270 ;
        RECT 2350.730 556.090 2351.910 557.270 ;
        RECT 2349.130 554.490 2350.310 555.670 ;
        RECT 2350.730 554.490 2351.910 555.670 ;
        RECT 2349.130 376.090 2350.310 377.270 ;
        RECT 2350.730 376.090 2351.910 377.270 ;
        RECT 2349.130 374.490 2350.310 375.670 ;
        RECT 2350.730 374.490 2351.910 375.670 ;
        RECT 2349.130 196.090 2350.310 197.270 ;
        RECT 2350.730 196.090 2351.910 197.270 ;
        RECT 2349.130 194.490 2350.310 195.670 ;
        RECT 2350.730 194.490 2351.910 195.670 ;
        RECT 2349.130 16.090 2350.310 17.270 ;
        RECT 2350.730 16.090 2351.910 17.270 ;
        RECT 2349.130 14.490 2350.310 15.670 ;
        RECT 2350.730 14.490 2351.910 15.670 ;
        RECT 2349.130 -2.910 2350.310 -1.730 ;
        RECT 2350.730 -2.910 2351.910 -1.730 ;
        RECT 2349.130 -4.510 2350.310 -3.330 ;
        RECT 2350.730 -4.510 2351.910 -3.330 ;
        RECT 2529.130 3523.010 2530.310 3524.190 ;
        RECT 2530.730 3523.010 2531.910 3524.190 ;
        RECT 2529.130 3521.410 2530.310 3522.590 ;
        RECT 2530.730 3521.410 2531.910 3522.590 ;
        RECT 2529.130 3436.090 2530.310 3437.270 ;
        RECT 2530.730 3436.090 2531.910 3437.270 ;
        RECT 2529.130 3434.490 2530.310 3435.670 ;
        RECT 2530.730 3434.490 2531.910 3435.670 ;
        RECT 2529.130 3256.090 2530.310 3257.270 ;
        RECT 2530.730 3256.090 2531.910 3257.270 ;
        RECT 2529.130 3254.490 2530.310 3255.670 ;
        RECT 2530.730 3254.490 2531.910 3255.670 ;
        RECT 2529.130 3076.090 2530.310 3077.270 ;
        RECT 2530.730 3076.090 2531.910 3077.270 ;
        RECT 2529.130 3074.490 2530.310 3075.670 ;
        RECT 2530.730 3074.490 2531.910 3075.670 ;
        RECT 2529.130 2896.090 2530.310 2897.270 ;
        RECT 2530.730 2896.090 2531.910 2897.270 ;
        RECT 2529.130 2894.490 2530.310 2895.670 ;
        RECT 2530.730 2894.490 2531.910 2895.670 ;
        RECT 2529.130 2716.090 2530.310 2717.270 ;
        RECT 2530.730 2716.090 2531.910 2717.270 ;
        RECT 2529.130 2714.490 2530.310 2715.670 ;
        RECT 2530.730 2714.490 2531.910 2715.670 ;
        RECT 2529.130 2536.090 2530.310 2537.270 ;
        RECT 2530.730 2536.090 2531.910 2537.270 ;
        RECT 2529.130 2534.490 2530.310 2535.670 ;
        RECT 2530.730 2534.490 2531.910 2535.670 ;
        RECT 2529.130 2356.090 2530.310 2357.270 ;
        RECT 2530.730 2356.090 2531.910 2357.270 ;
        RECT 2529.130 2354.490 2530.310 2355.670 ;
        RECT 2530.730 2354.490 2531.910 2355.670 ;
        RECT 2529.130 2176.090 2530.310 2177.270 ;
        RECT 2530.730 2176.090 2531.910 2177.270 ;
        RECT 2529.130 2174.490 2530.310 2175.670 ;
        RECT 2530.730 2174.490 2531.910 2175.670 ;
        RECT 2529.130 1996.090 2530.310 1997.270 ;
        RECT 2530.730 1996.090 2531.910 1997.270 ;
        RECT 2529.130 1994.490 2530.310 1995.670 ;
        RECT 2530.730 1994.490 2531.910 1995.670 ;
        RECT 2529.130 1816.090 2530.310 1817.270 ;
        RECT 2530.730 1816.090 2531.910 1817.270 ;
        RECT 2529.130 1814.490 2530.310 1815.670 ;
        RECT 2530.730 1814.490 2531.910 1815.670 ;
        RECT 2529.130 1636.090 2530.310 1637.270 ;
        RECT 2530.730 1636.090 2531.910 1637.270 ;
        RECT 2529.130 1634.490 2530.310 1635.670 ;
        RECT 2530.730 1634.490 2531.910 1635.670 ;
        RECT 2529.130 1456.090 2530.310 1457.270 ;
        RECT 2530.730 1456.090 2531.910 1457.270 ;
        RECT 2529.130 1454.490 2530.310 1455.670 ;
        RECT 2530.730 1454.490 2531.910 1455.670 ;
        RECT 2529.130 1276.090 2530.310 1277.270 ;
        RECT 2530.730 1276.090 2531.910 1277.270 ;
        RECT 2529.130 1274.490 2530.310 1275.670 ;
        RECT 2530.730 1274.490 2531.910 1275.670 ;
        RECT 2529.130 1096.090 2530.310 1097.270 ;
        RECT 2530.730 1096.090 2531.910 1097.270 ;
        RECT 2529.130 1094.490 2530.310 1095.670 ;
        RECT 2530.730 1094.490 2531.910 1095.670 ;
        RECT 2529.130 916.090 2530.310 917.270 ;
        RECT 2530.730 916.090 2531.910 917.270 ;
        RECT 2529.130 914.490 2530.310 915.670 ;
        RECT 2530.730 914.490 2531.910 915.670 ;
        RECT 2529.130 736.090 2530.310 737.270 ;
        RECT 2530.730 736.090 2531.910 737.270 ;
        RECT 2529.130 734.490 2530.310 735.670 ;
        RECT 2530.730 734.490 2531.910 735.670 ;
        RECT 2529.130 556.090 2530.310 557.270 ;
        RECT 2530.730 556.090 2531.910 557.270 ;
        RECT 2529.130 554.490 2530.310 555.670 ;
        RECT 2530.730 554.490 2531.910 555.670 ;
        RECT 2529.130 376.090 2530.310 377.270 ;
        RECT 2530.730 376.090 2531.910 377.270 ;
        RECT 2529.130 374.490 2530.310 375.670 ;
        RECT 2530.730 374.490 2531.910 375.670 ;
        RECT 2529.130 196.090 2530.310 197.270 ;
        RECT 2530.730 196.090 2531.910 197.270 ;
        RECT 2529.130 194.490 2530.310 195.670 ;
        RECT 2530.730 194.490 2531.910 195.670 ;
        RECT 2529.130 16.090 2530.310 17.270 ;
        RECT 2530.730 16.090 2531.910 17.270 ;
        RECT 2529.130 14.490 2530.310 15.670 ;
        RECT 2530.730 14.490 2531.910 15.670 ;
        RECT 2529.130 -2.910 2530.310 -1.730 ;
        RECT 2530.730 -2.910 2531.910 -1.730 ;
        RECT 2529.130 -4.510 2530.310 -3.330 ;
        RECT 2530.730 -4.510 2531.910 -3.330 ;
        RECT 2709.130 3523.010 2710.310 3524.190 ;
        RECT 2710.730 3523.010 2711.910 3524.190 ;
        RECT 2709.130 3521.410 2710.310 3522.590 ;
        RECT 2710.730 3521.410 2711.910 3522.590 ;
        RECT 2709.130 3436.090 2710.310 3437.270 ;
        RECT 2710.730 3436.090 2711.910 3437.270 ;
        RECT 2709.130 3434.490 2710.310 3435.670 ;
        RECT 2710.730 3434.490 2711.910 3435.670 ;
        RECT 2709.130 3256.090 2710.310 3257.270 ;
        RECT 2710.730 3256.090 2711.910 3257.270 ;
        RECT 2709.130 3254.490 2710.310 3255.670 ;
        RECT 2710.730 3254.490 2711.910 3255.670 ;
        RECT 2709.130 3076.090 2710.310 3077.270 ;
        RECT 2710.730 3076.090 2711.910 3077.270 ;
        RECT 2709.130 3074.490 2710.310 3075.670 ;
        RECT 2710.730 3074.490 2711.910 3075.670 ;
        RECT 2709.130 2896.090 2710.310 2897.270 ;
        RECT 2710.730 2896.090 2711.910 2897.270 ;
        RECT 2709.130 2894.490 2710.310 2895.670 ;
        RECT 2710.730 2894.490 2711.910 2895.670 ;
        RECT 2709.130 2716.090 2710.310 2717.270 ;
        RECT 2710.730 2716.090 2711.910 2717.270 ;
        RECT 2709.130 2714.490 2710.310 2715.670 ;
        RECT 2710.730 2714.490 2711.910 2715.670 ;
        RECT 2709.130 2536.090 2710.310 2537.270 ;
        RECT 2710.730 2536.090 2711.910 2537.270 ;
        RECT 2709.130 2534.490 2710.310 2535.670 ;
        RECT 2710.730 2534.490 2711.910 2535.670 ;
        RECT 2709.130 2356.090 2710.310 2357.270 ;
        RECT 2710.730 2356.090 2711.910 2357.270 ;
        RECT 2709.130 2354.490 2710.310 2355.670 ;
        RECT 2710.730 2354.490 2711.910 2355.670 ;
        RECT 2709.130 2176.090 2710.310 2177.270 ;
        RECT 2710.730 2176.090 2711.910 2177.270 ;
        RECT 2709.130 2174.490 2710.310 2175.670 ;
        RECT 2710.730 2174.490 2711.910 2175.670 ;
        RECT 2709.130 1996.090 2710.310 1997.270 ;
        RECT 2710.730 1996.090 2711.910 1997.270 ;
        RECT 2709.130 1994.490 2710.310 1995.670 ;
        RECT 2710.730 1994.490 2711.910 1995.670 ;
        RECT 2709.130 1816.090 2710.310 1817.270 ;
        RECT 2710.730 1816.090 2711.910 1817.270 ;
        RECT 2709.130 1814.490 2710.310 1815.670 ;
        RECT 2710.730 1814.490 2711.910 1815.670 ;
        RECT 2709.130 1636.090 2710.310 1637.270 ;
        RECT 2710.730 1636.090 2711.910 1637.270 ;
        RECT 2709.130 1634.490 2710.310 1635.670 ;
        RECT 2710.730 1634.490 2711.910 1635.670 ;
        RECT 2709.130 1456.090 2710.310 1457.270 ;
        RECT 2710.730 1456.090 2711.910 1457.270 ;
        RECT 2709.130 1454.490 2710.310 1455.670 ;
        RECT 2710.730 1454.490 2711.910 1455.670 ;
        RECT 2709.130 1276.090 2710.310 1277.270 ;
        RECT 2710.730 1276.090 2711.910 1277.270 ;
        RECT 2709.130 1274.490 2710.310 1275.670 ;
        RECT 2710.730 1274.490 2711.910 1275.670 ;
        RECT 2709.130 1096.090 2710.310 1097.270 ;
        RECT 2710.730 1096.090 2711.910 1097.270 ;
        RECT 2709.130 1094.490 2710.310 1095.670 ;
        RECT 2710.730 1094.490 2711.910 1095.670 ;
        RECT 2709.130 916.090 2710.310 917.270 ;
        RECT 2710.730 916.090 2711.910 917.270 ;
        RECT 2709.130 914.490 2710.310 915.670 ;
        RECT 2710.730 914.490 2711.910 915.670 ;
        RECT 2709.130 736.090 2710.310 737.270 ;
        RECT 2710.730 736.090 2711.910 737.270 ;
        RECT 2709.130 734.490 2710.310 735.670 ;
        RECT 2710.730 734.490 2711.910 735.670 ;
        RECT 2709.130 556.090 2710.310 557.270 ;
        RECT 2710.730 556.090 2711.910 557.270 ;
        RECT 2709.130 554.490 2710.310 555.670 ;
        RECT 2710.730 554.490 2711.910 555.670 ;
        RECT 2709.130 376.090 2710.310 377.270 ;
        RECT 2710.730 376.090 2711.910 377.270 ;
        RECT 2709.130 374.490 2710.310 375.670 ;
        RECT 2710.730 374.490 2711.910 375.670 ;
        RECT 2709.130 196.090 2710.310 197.270 ;
        RECT 2710.730 196.090 2711.910 197.270 ;
        RECT 2709.130 194.490 2710.310 195.670 ;
        RECT 2710.730 194.490 2711.910 195.670 ;
        RECT 2709.130 16.090 2710.310 17.270 ;
        RECT 2710.730 16.090 2711.910 17.270 ;
        RECT 2709.130 14.490 2710.310 15.670 ;
        RECT 2710.730 14.490 2711.910 15.670 ;
        RECT 2709.130 -2.910 2710.310 -1.730 ;
        RECT 2710.730 -2.910 2711.910 -1.730 ;
        RECT 2709.130 -4.510 2710.310 -3.330 ;
        RECT 2710.730 -4.510 2711.910 -3.330 ;
        RECT 2889.130 3523.010 2890.310 3524.190 ;
        RECT 2890.730 3523.010 2891.910 3524.190 ;
        RECT 2889.130 3521.410 2890.310 3522.590 ;
        RECT 2890.730 3521.410 2891.910 3522.590 ;
        RECT 2889.130 3436.090 2890.310 3437.270 ;
        RECT 2890.730 3436.090 2891.910 3437.270 ;
        RECT 2889.130 3434.490 2890.310 3435.670 ;
        RECT 2890.730 3434.490 2891.910 3435.670 ;
        RECT 2889.130 3256.090 2890.310 3257.270 ;
        RECT 2890.730 3256.090 2891.910 3257.270 ;
        RECT 2889.130 3254.490 2890.310 3255.670 ;
        RECT 2890.730 3254.490 2891.910 3255.670 ;
        RECT 2889.130 3076.090 2890.310 3077.270 ;
        RECT 2890.730 3076.090 2891.910 3077.270 ;
        RECT 2889.130 3074.490 2890.310 3075.670 ;
        RECT 2890.730 3074.490 2891.910 3075.670 ;
        RECT 2889.130 2896.090 2890.310 2897.270 ;
        RECT 2890.730 2896.090 2891.910 2897.270 ;
        RECT 2889.130 2894.490 2890.310 2895.670 ;
        RECT 2890.730 2894.490 2891.910 2895.670 ;
        RECT 2889.130 2716.090 2890.310 2717.270 ;
        RECT 2890.730 2716.090 2891.910 2717.270 ;
        RECT 2889.130 2714.490 2890.310 2715.670 ;
        RECT 2890.730 2714.490 2891.910 2715.670 ;
        RECT 2889.130 2536.090 2890.310 2537.270 ;
        RECT 2890.730 2536.090 2891.910 2537.270 ;
        RECT 2889.130 2534.490 2890.310 2535.670 ;
        RECT 2890.730 2534.490 2891.910 2535.670 ;
        RECT 2889.130 2356.090 2890.310 2357.270 ;
        RECT 2890.730 2356.090 2891.910 2357.270 ;
        RECT 2889.130 2354.490 2890.310 2355.670 ;
        RECT 2890.730 2354.490 2891.910 2355.670 ;
        RECT 2889.130 2176.090 2890.310 2177.270 ;
        RECT 2890.730 2176.090 2891.910 2177.270 ;
        RECT 2889.130 2174.490 2890.310 2175.670 ;
        RECT 2890.730 2174.490 2891.910 2175.670 ;
        RECT 2889.130 1996.090 2890.310 1997.270 ;
        RECT 2890.730 1996.090 2891.910 1997.270 ;
        RECT 2889.130 1994.490 2890.310 1995.670 ;
        RECT 2890.730 1994.490 2891.910 1995.670 ;
        RECT 2889.130 1816.090 2890.310 1817.270 ;
        RECT 2890.730 1816.090 2891.910 1817.270 ;
        RECT 2889.130 1814.490 2890.310 1815.670 ;
        RECT 2890.730 1814.490 2891.910 1815.670 ;
        RECT 2889.130 1636.090 2890.310 1637.270 ;
        RECT 2890.730 1636.090 2891.910 1637.270 ;
        RECT 2889.130 1634.490 2890.310 1635.670 ;
        RECT 2890.730 1634.490 2891.910 1635.670 ;
        RECT 2889.130 1456.090 2890.310 1457.270 ;
        RECT 2890.730 1456.090 2891.910 1457.270 ;
        RECT 2889.130 1454.490 2890.310 1455.670 ;
        RECT 2890.730 1454.490 2891.910 1455.670 ;
        RECT 2889.130 1276.090 2890.310 1277.270 ;
        RECT 2890.730 1276.090 2891.910 1277.270 ;
        RECT 2889.130 1274.490 2890.310 1275.670 ;
        RECT 2890.730 1274.490 2891.910 1275.670 ;
        RECT 2889.130 1096.090 2890.310 1097.270 ;
        RECT 2890.730 1096.090 2891.910 1097.270 ;
        RECT 2889.130 1094.490 2890.310 1095.670 ;
        RECT 2890.730 1094.490 2891.910 1095.670 ;
        RECT 2889.130 916.090 2890.310 917.270 ;
        RECT 2890.730 916.090 2891.910 917.270 ;
        RECT 2889.130 914.490 2890.310 915.670 ;
        RECT 2890.730 914.490 2891.910 915.670 ;
        RECT 2889.130 736.090 2890.310 737.270 ;
        RECT 2890.730 736.090 2891.910 737.270 ;
        RECT 2889.130 734.490 2890.310 735.670 ;
        RECT 2890.730 734.490 2891.910 735.670 ;
        RECT 2889.130 556.090 2890.310 557.270 ;
        RECT 2890.730 556.090 2891.910 557.270 ;
        RECT 2889.130 554.490 2890.310 555.670 ;
        RECT 2890.730 554.490 2891.910 555.670 ;
        RECT 2889.130 376.090 2890.310 377.270 ;
        RECT 2890.730 376.090 2891.910 377.270 ;
        RECT 2889.130 374.490 2890.310 375.670 ;
        RECT 2890.730 374.490 2891.910 375.670 ;
        RECT 2889.130 196.090 2890.310 197.270 ;
        RECT 2890.730 196.090 2891.910 197.270 ;
        RECT 2889.130 194.490 2890.310 195.670 ;
        RECT 2890.730 194.490 2891.910 195.670 ;
        RECT 2889.130 16.090 2890.310 17.270 ;
        RECT 2890.730 16.090 2891.910 17.270 ;
        RECT 2889.130 14.490 2890.310 15.670 ;
        RECT 2890.730 14.490 2891.910 15.670 ;
        RECT 2889.130 -2.910 2890.310 -1.730 ;
        RECT 2890.730 -2.910 2891.910 -1.730 ;
        RECT 2889.130 -4.510 2890.310 -3.330 ;
        RECT 2890.730 -4.510 2891.910 -3.330 ;
        RECT 2926.710 3523.010 2927.890 3524.190 ;
        RECT 2928.310 3523.010 2929.490 3524.190 ;
        RECT 2926.710 3521.410 2927.890 3522.590 ;
        RECT 2928.310 3521.410 2929.490 3522.590 ;
        RECT 2926.710 3436.090 2927.890 3437.270 ;
        RECT 2928.310 3436.090 2929.490 3437.270 ;
        RECT 2926.710 3434.490 2927.890 3435.670 ;
        RECT 2928.310 3434.490 2929.490 3435.670 ;
        RECT 2926.710 3256.090 2927.890 3257.270 ;
        RECT 2928.310 3256.090 2929.490 3257.270 ;
        RECT 2926.710 3254.490 2927.890 3255.670 ;
        RECT 2928.310 3254.490 2929.490 3255.670 ;
        RECT 2926.710 3076.090 2927.890 3077.270 ;
        RECT 2928.310 3076.090 2929.490 3077.270 ;
        RECT 2926.710 3074.490 2927.890 3075.670 ;
        RECT 2928.310 3074.490 2929.490 3075.670 ;
        RECT 2926.710 2896.090 2927.890 2897.270 ;
        RECT 2928.310 2896.090 2929.490 2897.270 ;
        RECT 2926.710 2894.490 2927.890 2895.670 ;
        RECT 2928.310 2894.490 2929.490 2895.670 ;
        RECT 2926.710 2716.090 2927.890 2717.270 ;
        RECT 2928.310 2716.090 2929.490 2717.270 ;
        RECT 2926.710 2714.490 2927.890 2715.670 ;
        RECT 2928.310 2714.490 2929.490 2715.670 ;
        RECT 2926.710 2536.090 2927.890 2537.270 ;
        RECT 2928.310 2536.090 2929.490 2537.270 ;
        RECT 2926.710 2534.490 2927.890 2535.670 ;
        RECT 2928.310 2534.490 2929.490 2535.670 ;
        RECT 2926.710 2356.090 2927.890 2357.270 ;
        RECT 2928.310 2356.090 2929.490 2357.270 ;
        RECT 2926.710 2354.490 2927.890 2355.670 ;
        RECT 2928.310 2354.490 2929.490 2355.670 ;
        RECT 2926.710 2176.090 2927.890 2177.270 ;
        RECT 2928.310 2176.090 2929.490 2177.270 ;
        RECT 2926.710 2174.490 2927.890 2175.670 ;
        RECT 2928.310 2174.490 2929.490 2175.670 ;
        RECT 2926.710 1996.090 2927.890 1997.270 ;
        RECT 2928.310 1996.090 2929.490 1997.270 ;
        RECT 2926.710 1994.490 2927.890 1995.670 ;
        RECT 2928.310 1994.490 2929.490 1995.670 ;
        RECT 2926.710 1816.090 2927.890 1817.270 ;
        RECT 2928.310 1816.090 2929.490 1817.270 ;
        RECT 2926.710 1814.490 2927.890 1815.670 ;
        RECT 2928.310 1814.490 2929.490 1815.670 ;
        RECT 2926.710 1636.090 2927.890 1637.270 ;
        RECT 2928.310 1636.090 2929.490 1637.270 ;
        RECT 2926.710 1634.490 2927.890 1635.670 ;
        RECT 2928.310 1634.490 2929.490 1635.670 ;
        RECT 2926.710 1456.090 2927.890 1457.270 ;
        RECT 2928.310 1456.090 2929.490 1457.270 ;
        RECT 2926.710 1454.490 2927.890 1455.670 ;
        RECT 2928.310 1454.490 2929.490 1455.670 ;
        RECT 2926.710 1276.090 2927.890 1277.270 ;
        RECT 2928.310 1276.090 2929.490 1277.270 ;
        RECT 2926.710 1274.490 2927.890 1275.670 ;
        RECT 2928.310 1274.490 2929.490 1275.670 ;
        RECT 2926.710 1096.090 2927.890 1097.270 ;
        RECT 2928.310 1096.090 2929.490 1097.270 ;
        RECT 2926.710 1094.490 2927.890 1095.670 ;
        RECT 2928.310 1094.490 2929.490 1095.670 ;
        RECT 2926.710 916.090 2927.890 917.270 ;
        RECT 2928.310 916.090 2929.490 917.270 ;
        RECT 2926.710 914.490 2927.890 915.670 ;
        RECT 2928.310 914.490 2929.490 915.670 ;
        RECT 2926.710 736.090 2927.890 737.270 ;
        RECT 2928.310 736.090 2929.490 737.270 ;
        RECT 2926.710 734.490 2927.890 735.670 ;
        RECT 2928.310 734.490 2929.490 735.670 ;
        RECT 2926.710 556.090 2927.890 557.270 ;
        RECT 2928.310 556.090 2929.490 557.270 ;
        RECT 2926.710 554.490 2927.890 555.670 ;
        RECT 2928.310 554.490 2929.490 555.670 ;
        RECT 2926.710 376.090 2927.890 377.270 ;
        RECT 2928.310 376.090 2929.490 377.270 ;
        RECT 2926.710 374.490 2927.890 375.670 ;
        RECT 2928.310 374.490 2929.490 375.670 ;
        RECT 2926.710 196.090 2927.890 197.270 ;
        RECT 2928.310 196.090 2929.490 197.270 ;
        RECT 2926.710 194.490 2927.890 195.670 ;
        RECT 2928.310 194.490 2929.490 195.670 ;
        RECT 2926.710 16.090 2927.890 17.270 ;
        RECT 2928.310 16.090 2929.490 17.270 ;
        RECT 2926.710 14.490 2927.890 15.670 ;
        RECT 2928.310 14.490 2929.490 15.670 ;
        RECT 2926.710 -2.910 2927.890 -1.730 ;
        RECT 2928.310 -2.910 2929.490 -1.730 ;
        RECT 2926.710 -4.510 2927.890 -3.330 ;
        RECT 2928.310 -4.510 2929.490 -3.330 ;
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
        RECT -43.630 3434.330 2963.250 3437.430 ;
        RECT -43.630 3254.330 2963.250 3257.430 ;
        RECT -43.630 3074.330 2963.250 3077.430 ;
        RECT -43.630 2894.330 2963.250 2897.430 ;
        RECT -43.630 2714.330 2963.250 2717.430 ;
        RECT -43.630 2534.330 2963.250 2537.430 ;
        RECT -43.630 2354.330 2963.250 2357.430 ;
        RECT -43.630 2174.330 2963.250 2177.430 ;
        RECT -43.630 1994.330 2963.250 1997.430 ;
        RECT -43.630 1814.330 2963.250 1817.430 ;
        RECT -43.630 1634.330 2963.250 1637.430 ;
        RECT -43.630 1454.330 2963.250 1457.430 ;
        RECT -43.630 1274.330 2963.250 1277.430 ;
        RECT -43.630 1094.330 2963.250 1097.430 ;
        RECT -43.630 914.330 2963.250 917.430 ;
        RECT -43.630 734.330 2963.250 737.430 ;
        RECT -43.630 554.330 2963.250 557.430 ;
        RECT -43.630 374.330 2963.250 377.430 ;
        RECT -43.630 194.330 2963.250 197.430 ;
        RECT -43.630 14.330 2963.250 17.430 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
        RECT 53.970 -38.270 57.070 3557.950 ;
        RECT 233.970 -38.270 237.070 3557.950 ;
        RECT 413.970 810.000 417.070 3557.950 ;
        RECT 593.970 810.000 597.070 3557.950 ;
        RECT 413.970 -38.270 417.070 490.000 ;
        RECT 593.970 -38.270 597.070 490.000 ;
        RECT 773.970 -38.270 777.070 3557.950 ;
        RECT 953.970 -38.270 957.070 3557.950 ;
        RECT 1133.970 -38.270 1137.070 3557.950 ;
        RECT 1313.970 -38.270 1317.070 3557.950 ;
        RECT 1493.970 -38.270 1497.070 3557.950 ;
        RECT 1673.970 -38.270 1677.070 3557.950 ;
        RECT 1853.970 -38.270 1857.070 3557.950 ;
        RECT 2033.970 -38.270 2037.070 3557.950 ;
        RECT 2213.970 -38.270 2217.070 3557.950 ;
        RECT 2393.970 -38.270 2397.070 3557.950 ;
        RECT 2573.970 -38.270 2577.070 3557.950 ;
        RECT 2753.970 -38.270 2757.070 3557.950 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
      LAYER via4 ;
        RECT -19.470 3532.610 -18.290 3533.790 ;
        RECT -17.870 3532.610 -16.690 3533.790 ;
        RECT -19.470 3531.010 -18.290 3532.190 ;
        RECT -17.870 3531.010 -16.690 3532.190 ;
        RECT -19.470 3481.090 -18.290 3482.270 ;
        RECT -17.870 3481.090 -16.690 3482.270 ;
        RECT -19.470 3479.490 -18.290 3480.670 ;
        RECT -17.870 3479.490 -16.690 3480.670 ;
        RECT -19.470 3301.090 -18.290 3302.270 ;
        RECT -17.870 3301.090 -16.690 3302.270 ;
        RECT -19.470 3299.490 -18.290 3300.670 ;
        RECT -17.870 3299.490 -16.690 3300.670 ;
        RECT -19.470 3121.090 -18.290 3122.270 ;
        RECT -17.870 3121.090 -16.690 3122.270 ;
        RECT -19.470 3119.490 -18.290 3120.670 ;
        RECT -17.870 3119.490 -16.690 3120.670 ;
        RECT -19.470 2941.090 -18.290 2942.270 ;
        RECT -17.870 2941.090 -16.690 2942.270 ;
        RECT -19.470 2939.490 -18.290 2940.670 ;
        RECT -17.870 2939.490 -16.690 2940.670 ;
        RECT -19.470 2761.090 -18.290 2762.270 ;
        RECT -17.870 2761.090 -16.690 2762.270 ;
        RECT -19.470 2759.490 -18.290 2760.670 ;
        RECT -17.870 2759.490 -16.690 2760.670 ;
        RECT -19.470 2581.090 -18.290 2582.270 ;
        RECT -17.870 2581.090 -16.690 2582.270 ;
        RECT -19.470 2579.490 -18.290 2580.670 ;
        RECT -17.870 2579.490 -16.690 2580.670 ;
        RECT -19.470 2401.090 -18.290 2402.270 ;
        RECT -17.870 2401.090 -16.690 2402.270 ;
        RECT -19.470 2399.490 -18.290 2400.670 ;
        RECT -17.870 2399.490 -16.690 2400.670 ;
        RECT -19.470 2221.090 -18.290 2222.270 ;
        RECT -17.870 2221.090 -16.690 2222.270 ;
        RECT -19.470 2219.490 -18.290 2220.670 ;
        RECT -17.870 2219.490 -16.690 2220.670 ;
        RECT -19.470 2041.090 -18.290 2042.270 ;
        RECT -17.870 2041.090 -16.690 2042.270 ;
        RECT -19.470 2039.490 -18.290 2040.670 ;
        RECT -17.870 2039.490 -16.690 2040.670 ;
        RECT -19.470 1861.090 -18.290 1862.270 ;
        RECT -17.870 1861.090 -16.690 1862.270 ;
        RECT -19.470 1859.490 -18.290 1860.670 ;
        RECT -17.870 1859.490 -16.690 1860.670 ;
        RECT -19.470 1681.090 -18.290 1682.270 ;
        RECT -17.870 1681.090 -16.690 1682.270 ;
        RECT -19.470 1679.490 -18.290 1680.670 ;
        RECT -17.870 1679.490 -16.690 1680.670 ;
        RECT -19.470 1501.090 -18.290 1502.270 ;
        RECT -17.870 1501.090 -16.690 1502.270 ;
        RECT -19.470 1499.490 -18.290 1500.670 ;
        RECT -17.870 1499.490 -16.690 1500.670 ;
        RECT -19.470 1321.090 -18.290 1322.270 ;
        RECT -17.870 1321.090 -16.690 1322.270 ;
        RECT -19.470 1319.490 -18.290 1320.670 ;
        RECT -17.870 1319.490 -16.690 1320.670 ;
        RECT -19.470 1141.090 -18.290 1142.270 ;
        RECT -17.870 1141.090 -16.690 1142.270 ;
        RECT -19.470 1139.490 -18.290 1140.670 ;
        RECT -17.870 1139.490 -16.690 1140.670 ;
        RECT -19.470 961.090 -18.290 962.270 ;
        RECT -17.870 961.090 -16.690 962.270 ;
        RECT -19.470 959.490 -18.290 960.670 ;
        RECT -17.870 959.490 -16.690 960.670 ;
        RECT -19.470 781.090 -18.290 782.270 ;
        RECT -17.870 781.090 -16.690 782.270 ;
        RECT -19.470 779.490 -18.290 780.670 ;
        RECT -17.870 779.490 -16.690 780.670 ;
        RECT -19.470 601.090 -18.290 602.270 ;
        RECT -17.870 601.090 -16.690 602.270 ;
        RECT -19.470 599.490 -18.290 600.670 ;
        RECT -17.870 599.490 -16.690 600.670 ;
        RECT -19.470 421.090 -18.290 422.270 ;
        RECT -17.870 421.090 -16.690 422.270 ;
        RECT -19.470 419.490 -18.290 420.670 ;
        RECT -17.870 419.490 -16.690 420.670 ;
        RECT -19.470 241.090 -18.290 242.270 ;
        RECT -17.870 241.090 -16.690 242.270 ;
        RECT -19.470 239.490 -18.290 240.670 ;
        RECT -17.870 239.490 -16.690 240.670 ;
        RECT -19.470 61.090 -18.290 62.270 ;
        RECT -17.870 61.090 -16.690 62.270 ;
        RECT -19.470 59.490 -18.290 60.670 ;
        RECT -17.870 59.490 -16.690 60.670 ;
        RECT -19.470 -12.510 -18.290 -11.330 ;
        RECT -17.870 -12.510 -16.690 -11.330 ;
        RECT -19.470 -14.110 -18.290 -12.930 ;
        RECT -17.870 -14.110 -16.690 -12.930 ;
        RECT 54.130 3532.610 55.310 3533.790 ;
        RECT 55.730 3532.610 56.910 3533.790 ;
        RECT 54.130 3531.010 55.310 3532.190 ;
        RECT 55.730 3531.010 56.910 3532.190 ;
        RECT 54.130 3481.090 55.310 3482.270 ;
        RECT 55.730 3481.090 56.910 3482.270 ;
        RECT 54.130 3479.490 55.310 3480.670 ;
        RECT 55.730 3479.490 56.910 3480.670 ;
        RECT 54.130 3301.090 55.310 3302.270 ;
        RECT 55.730 3301.090 56.910 3302.270 ;
        RECT 54.130 3299.490 55.310 3300.670 ;
        RECT 55.730 3299.490 56.910 3300.670 ;
        RECT 54.130 3121.090 55.310 3122.270 ;
        RECT 55.730 3121.090 56.910 3122.270 ;
        RECT 54.130 3119.490 55.310 3120.670 ;
        RECT 55.730 3119.490 56.910 3120.670 ;
        RECT 54.130 2941.090 55.310 2942.270 ;
        RECT 55.730 2941.090 56.910 2942.270 ;
        RECT 54.130 2939.490 55.310 2940.670 ;
        RECT 55.730 2939.490 56.910 2940.670 ;
        RECT 54.130 2761.090 55.310 2762.270 ;
        RECT 55.730 2761.090 56.910 2762.270 ;
        RECT 54.130 2759.490 55.310 2760.670 ;
        RECT 55.730 2759.490 56.910 2760.670 ;
        RECT 54.130 2581.090 55.310 2582.270 ;
        RECT 55.730 2581.090 56.910 2582.270 ;
        RECT 54.130 2579.490 55.310 2580.670 ;
        RECT 55.730 2579.490 56.910 2580.670 ;
        RECT 54.130 2401.090 55.310 2402.270 ;
        RECT 55.730 2401.090 56.910 2402.270 ;
        RECT 54.130 2399.490 55.310 2400.670 ;
        RECT 55.730 2399.490 56.910 2400.670 ;
        RECT 54.130 2221.090 55.310 2222.270 ;
        RECT 55.730 2221.090 56.910 2222.270 ;
        RECT 54.130 2219.490 55.310 2220.670 ;
        RECT 55.730 2219.490 56.910 2220.670 ;
        RECT 54.130 2041.090 55.310 2042.270 ;
        RECT 55.730 2041.090 56.910 2042.270 ;
        RECT 54.130 2039.490 55.310 2040.670 ;
        RECT 55.730 2039.490 56.910 2040.670 ;
        RECT 54.130 1861.090 55.310 1862.270 ;
        RECT 55.730 1861.090 56.910 1862.270 ;
        RECT 54.130 1859.490 55.310 1860.670 ;
        RECT 55.730 1859.490 56.910 1860.670 ;
        RECT 54.130 1681.090 55.310 1682.270 ;
        RECT 55.730 1681.090 56.910 1682.270 ;
        RECT 54.130 1679.490 55.310 1680.670 ;
        RECT 55.730 1679.490 56.910 1680.670 ;
        RECT 54.130 1501.090 55.310 1502.270 ;
        RECT 55.730 1501.090 56.910 1502.270 ;
        RECT 54.130 1499.490 55.310 1500.670 ;
        RECT 55.730 1499.490 56.910 1500.670 ;
        RECT 54.130 1321.090 55.310 1322.270 ;
        RECT 55.730 1321.090 56.910 1322.270 ;
        RECT 54.130 1319.490 55.310 1320.670 ;
        RECT 55.730 1319.490 56.910 1320.670 ;
        RECT 54.130 1141.090 55.310 1142.270 ;
        RECT 55.730 1141.090 56.910 1142.270 ;
        RECT 54.130 1139.490 55.310 1140.670 ;
        RECT 55.730 1139.490 56.910 1140.670 ;
        RECT 54.130 961.090 55.310 962.270 ;
        RECT 55.730 961.090 56.910 962.270 ;
        RECT 54.130 959.490 55.310 960.670 ;
        RECT 55.730 959.490 56.910 960.670 ;
        RECT 54.130 781.090 55.310 782.270 ;
        RECT 55.730 781.090 56.910 782.270 ;
        RECT 54.130 779.490 55.310 780.670 ;
        RECT 55.730 779.490 56.910 780.670 ;
        RECT 54.130 601.090 55.310 602.270 ;
        RECT 55.730 601.090 56.910 602.270 ;
        RECT 54.130 599.490 55.310 600.670 ;
        RECT 55.730 599.490 56.910 600.670 ;
        RECT 54.130 421.090 55.310 422.270 ;
        RECT 55.730 421.090 56.910 422.270 ;
        RECT 54.130 419.490 55.310 420.670 ;
        RECT 55.730 419.490 56.910 420.670 ;
        RECT 54.130 241.090 55.310 242.270 ;
        RECT 55.730 241.090 56.910 242.270 ;
        RECT 54.130 239.490 55.310 240.670 ;
        RECT 55.730 239.490 56.910 240.670 ;
        RECT 54.130 61.090 55.310 62.270 ;
        RECT 55.730 61.090 56.910 62.270 ;
        RECT 54.130 59.490 55.310 60.670 ;
        RECT 55.730 59.490 56.910 60.670 ;
        RECT 54.130 -12.510 55.310 -11.330 ;
        RECT 55.730 -12.510 56.910 -11.330 ;
        RECT 54.130 -14.110 55.310 -12.930 ;
        RECT 55.730 -14.110 56.910 -12.930 ;
        RECT 234.130 3532.610 235.310 3533.790 ;
        RECT 235.730 3532.610 236.910 3533.790 ;
        RECT 234.130 3531.010 235.310 3532.190 ;
        RECT 235.730 3531.010 236.910 3532.190 ;
        RECT 234.130 3481.090 235.310 3482.270 ;
        RECT 235.730 3481.090 236.910 3482.270 ;
        RECT 234.130 3479.490 235.310 3480.670 ;
        RECT 235.730 3479.490 236.910 3480.670 ;
        RECT 234.130 3301.090 235.310 3302.270 ;
        RECT 235.730 3301.090 236.910 3302.270 ;
        RECT 234.130 3299.490 235.310 3300.670 ;
        RECT 235.730 3299.490 236.910 3300.670 ;
        RECT 234.130 3121.090 235.310 3122.270 ;
        RECT 235.730 3121.090 236.910 3122.270 ;
        RECT 234.130 3119.490 235.310 3120.670 ;
        RECT 235.730 3119.490 236.910 3120.670 ;
        RECT 234.130 2941.090 235.310 2942.270 ;
        RECT 235.730 2941.090 236.910 2942.270 ;
        RECT 234.130 2939.490 235.310 2940.670 ;
        RECT 235.730 2939.490 236.910 2940.670 ;
        RECT 234.130 2761.090 235.310 2762.270 ;
        RECT 235.730 2761.090 236.910 2762.270 ;
        RECT 234.130 2759.490 235.310 2760.670 ;
        RECT 235.730 2759.490 236.910 2760.670 ;
        RECT 234.130 2581.090 235.310 2582.270 ;
        RECT 235.730 2581.090 236.910 2582.270 ;
        RECT 234.130 2579.490 235.310 2580.670 ;
        RECT 235.730 2579.490 236.910 2580.670 ;
        RECT 234.130 2401.090 235.310 2402.270 ;
        RECT 235.730 2401.090 236.910 2402.270 ;
        RECT 234.130 2399.490 235.310 2400.670 ;
        RECT 235.730 2399.490 236.910 2400.670 ;
        RECT 234.130 2221.090 235.310 2222.270 ;
        RECT 235.730 2221.090 236.910 2222.270 ;
        RECT 234.130 2219.490 235.310 2220.670 ;
        RECT 235.730 2219.490 236.910 2220.670 ;
        RECT 234.130 2041.090 235.310 2042.270 ;
        RECT 235.730 2041.090 236.910 2042.270 ;
        RECT 234.130 2039.490 235.310 2040.670 ;
        RECT 235.730 2039.490 236.910 2040.670 ;
        RECT 234.130 1861.090 235.310 1862.270 ;
        RECT 235.730 1861.090 236.910 1862.270 ;
        RECT 234.130 1859.490 235.310 1860.670 ;
        RECT 235.730 1859.490 236.910 1860.670 ;
        RECT 234.130 1681.090 235.310 1682.270 ;
        RECT 235.730 1681.090 236.910 1682.270 ;
        RECT 234.130 1679.490 235.310 1680.670 ;
        RECT 235.730 1679.490 236.910 1680.670 ;
        RECT 234.130 1501.090 235.310 1502.270 ;
        RECT 235.730 1501.090 236.910 1502.270 ;
        RECT 234.130 1499.490 235.310 1500.670 ;
        RECT 235.730 1499.490 236.910 1500.670 ;
        RECT 234.130 1321.090 235.310 1322.270 ;
        RECT 235.730 1321.090 236.910 1322.270 ;
        RECT 234.130 1319.490 235.310 1320.670 ;
        RECT 235.730 1319.490 236.910 1320.670 ;
        RECT 234.130 1141.090 235.310 1142.270 ;
        RECT 235.730 1141.090 236.910 1142.270 ;
        RECT 234.130 1139.490 235.310 1140.670 ;
        RECT 235.730 1139.490 236.910 1140.670 ;
        RECT 234.130 961.090 235.310 962.270 ;
        RECT 235.730 961.090 236.910 962.270 ;
        RECT 234.130 959.490 235.310 960.670 ;
        RECT 235.730 959.490 236.910 960.670 ;
        RECT 414.130 3532.610 415.310 3533.790 ;
        RECT 415.730 3532.610 416.910 3533.790 ;
        RECT 414.130 3531.010 415.310 3532.190 ;
        RECT 415.730 3531.010 416.910 3532.190 ;
        RECT 414.130 3481.090 415.310 3482.270 ;
        RECT 415.730 3481.090 416.910 3482.270 ;
        RECT 414.130 3479.490 415.310 3480.670 ;
        RECT 415.730 3479.490 416.910 3480.670 ;
        RECT 414.130 3301.090 415.310 3302.270 ;
        RECT 415.730 3301.090 416.910 3302.270 ;
        RECT 414.130 3299.490 415.310 3300.670 ;
        RECT 415.730 3299.490 416.910 3300.670 ;
        RECT 414.130 3121.090 415.310 3122.270 ;
        RECT 415.730 3121.090 416.910 3122.270 ;
        RECT 414.130 3119.490 415.310 3120.670 ;
        RECT 415.730 3119.490 416.910 3120.670 ;
        RECT 414.130 2941.090 415.310 2942.270 ;
        RECT 415.730 2941.090 416.910 2942.270 ;
        RECT 414.130 2939.490 415.310 2940.670 ;
        RECT 415.730 2939.490 416.910 2940.670 ;
        RECT 414.130 2761.090 415.310 2762.270 ;
        RECT 415.730 2761.090 416.910 2762.270 ;
        RECT 414.130 2759.490 415.310 2760.670 ;
        RECT 415.730 2759.490 416.910 2760.670 ;
        RECT 414.130 2581.090 415.310 2582.270 ;
        RECT 415.730 2581.090 416.910 2582.270 ;
        RECT 414.130 2579.490 415.310 2580.670 ;
        RECT 415.730 2579.490 416.910 2580.670 ;
        RECT 414.130 2401.090 415.310 2402.270 ;
        RECT 415.730 2401.090 416.910 2402.270 ;
        RECT 414.130 2399.490 415.310 2400.670 ;
        RECT 415.730 2399.490 416.910 2400.670 ;
        RECT 414.130 2221.090 415.310 2222.270 ;
        RECT 415.730 2221.090 416.910 2222.270 ;
        RECT 414.130 2219.490 415.310 2220.670 ;
        RECT 415.730 2219.490 416.910 2220.670 ;
        RECT 414.130 2041.090 415.310 2042.270 ;
        RECT 415.730 2041.090 416.910 2042.270 ;
        RECT 414.130 2039.490 415.310 2040.670 ;
        RECT 415.730 2039.490 416.910 2040.670 ;
        RECT 414.130 1861.090 415.310 1862.270 ;
        RECT 415.730 1861.090 416.910 1862.270 ;
        RECT 414.130 1859.490 415.310 1860.670 ;
        RECT 415.730 1859.490 416.910 1860.670 ;
        RECT 414.130 1681.090 415.310 1682.270 ;
        RECT 415.730 1681.090 416.910 1682.270 ;
        RECT 414.130 1679.490 415.310 1680.670 ;
        RECT 415.730 1679.490 416.910 1680.670 ;
        RECT 414.130 1501.090 415.310 1502.270 ;
        RECT 415.730 1501.090 416.910 1502.270 ;
        RECT 414.130 1499.490 415.310 1500.670 ;
        RECT 415.730 1499.490 416.910 1500.670 ;
        RECT 414.130 1321.090 415.310 1322.270 ;
        RECT 415.730 1321.090 416.910 1322.270 ;
        RECT 414.130 1319.490 415.310 1320.670 ;
        RECT 415.730 1319.490 416.910 1320.670 ;
        RECT 414.130 1141.090 415.310 1142.270 ;
        RECT 415.730 1141.090 416.910 1142.270 ;
        RECT 414.130 1139.490 415.310 1140.670 ;
        RECT 415.730 1139.490 416.910 1140.670 ;
        RECT 414.130 961.090 415.310 962.270 ;
        RECT 415.730 961.090 416.910 962.270 ;
        RECT 414.130 959.490 415.310 960.670 ;
        RECT 415.730 959.490 416.910 960.670 ;
        RECT 594.130 3532.610 595.310 3533.790 ;
        RECT 595.730 3532.610 596.910 3533.790 ;
        RECT 594.130 3531.010 595.310 3532.190 ;
        RECT 595.730 3531.010 596.910 3532.190 ;
        RECT 594.130 3481.090 595.310 3482.270 ;
        RECT 595.730 3481.090 596.910 3482.270 ;
        RECT 594.130 3479.490 595.310 3480.670 ;
        RECT 595.730 3479.490 596.910 3480.670 ;
        RECT 594.130 3301.090 595.310 3302.270 ;
        RECT 595.730 3301.090 596.910 3302.270 ;
        RECT 594.130 3299.490 595.310 3300.670 ;
        RECT 595.730 3299.490 596.910 3300.670 ;
        RECT 594.130 3121.090 595.310 3122.270 ;
        RECT 595.730 3121.090 596.910 3122.270 ;
        RECT 594.130 3119.490 595.310 3120.670 ;
        RECT 595.730 3119.490 596.910 3120.670 ;
        RECT 594.130 2941.090 595.310 2942.270 ;
        RECT 595.730 2941.090 596.910 2942.270 ;
        RECT 594.130 2939.490 595.310 2940.670 ;
        RECT 595.730 2939.490 596.910 2940.670 ;
        RECT 594.130 2761.090 595.310 2762.270 ;
        RECT 595.730 2761.090 596.910 2762.270 ;
        RECT 594.130 2759.490 595.310 2760.670 ;
        RECT 595.730 2759.490 596.910 2760.670 ;
        RECT 594.130 2581.090 595.310 2582.270 ;
        RECT 595.730 2581.090 596.910 2582.270 ;
        RECT 594.130 2579.490 595.310 2580.670 ;
        RECT 595.730 2579.490 596.910 2580.670 ;
        RECT 594.130 2401.090 595.310 2402.270 ;
        RECT 595.730 2401.090 596.910 2402.270 ;
        RECT 594.130 2399.490 595.310 2400.670 ;
        RECT 595.730 2399.490 596.910 2400.670 ;
        RECT 594.130 2221.090 595.310 2222.270 ;
        RECT 595.730 2221.090 596.910 2222.270 ;
        RECT 594.130 2219.490 595.310 2220.670 ;
        RECT 595.730 2219.490 596.910 2220.670 ;
        RECT 594.130 2041.090 595.310 2042.270 ;
        RECT 595.730 2041.090 596.910 2042.270 ;
        RECT 594.130 2039.490 595.310 2040.670 ;
        RECT 595.730 2039.490 596.910 2040.670 ;
        RECT 594.130 1861.090 595.310 1862.270 ;
        RECT 595.730 1861.090 596.910 1862.270 ;
        RECT 594.130 1859.490 595.310 1860.670 ;
        RECT 595.730 1859.490 596.910 1860.670 ;
        RECT 594.130 1681.090 595.310 1682.270 ;
        RECT 595.730 1681.090 596.910 1682.270 ;
        RECT 594.130 1679.490 595.310 1680.670 ;
        RECT 595.730 1679.490 596.910 1680.670 ;
        RECT 594.130 1501.090 595.310 1502.270 ;
        RECT 595.730 1501.090 596.910 1502.270 ;
        RECT 594.130 1499.490 595.310 1500.670 ;
        RECT 595.730 1499.490 596.910 1500.670 ;
        RECT 594.130 1321.090 595.310 1322.270 ;
        RECT 595.730 1321.090 596.910 1322.270 ;
        RECT 594.130 1319.490 595.310 1320.670 ;
        RECT 595.730 1319.490 596.910 1320.670 ;
        RECT 594.130 1141.090 595.310 1142.270 ;
        RECT 595.730 1141.090 596.910 1142.270 ;
        RECT 594.130 1139.490 595.310 1140.670 ;
        RECT 595.730 1139.490 596.910 1140.670 ;
        RECT 594.130 961.090 595.310 962.270 ;
        RECT 595.730 961.090 596.910 962.270 ;
        RECT 594.130 959.490 595.310 960.670 ;
        RECT 595.730 959.490 596.910 960.670 ;
        RECT 774.130 3532.610 775.310 3533.790 ;
        RECT 775.730 3532.610 776.910 3533.790 ;
        RECT 774.130 3531.010 775.310 3532.190 ;
        RECT 775.730 3531.010 776.910 3532.190 ;
        RECT 774.130 3481.090 775.310 3482.270 ;
        RECT 775.730 3481.090 776.910 3482.270 ;
        RECT 774.130 3479.490 775.310 3480.670 ;
        RECT 775.730 3479.490 776.910 3480.670 ;
        RECT 774.130 3301.090 775.310 3302.270 ;
        RECT 775.730 3301.090 776.910 3302.270 ;
        RECT 774.130 3299.490 775.310 3300.670 ;
        RECT 775.730 3299.490 776.910 3300.670 ;
        RECT 774.130 3121.090 775.310 3122.270 ;
        RECT 775.730 3121.090 776.910 3122.270 ;
        RECT 774.130 3119.490 775.310 3120.670 ;
        RECT 775.730 3119.490 776.910 3120.670 ;
        RECT 774.130 2941.090 775.310 2942.270 ;
        RECT 775.730 2941.090 776.910 2942.270 ;
        RECT 774.130 2939.490 775.310 2940.670 ;
        RECT 775.730 2939.490 776.910 2940.670 ;
        RECT 774.130 2761.090 775.310 2762.270 ;
        RECT 775.730 2761.090 776.910 2762.270 ;
        RECT 774.130 2759.490 775.310 2760.670 ;
        RECT 775.730 2759.490 776.910 2760.670 ;
        RECT 774.130 2581.090 775.310 2582.270 ;
        RECT 775.730 2581.090 776.910 2582.270 ;
        RECT 774.130 2579.490 775.310 2580.670 ;
        RECT 775.730 2579.490 776.910 2580.670 ;
        RECT 774.130 2401.090 775.310 2402.270 ;
        RECT 775.730 2401.090 776.910 2402.270 ;
        RECT 774.130 2399.490 775.310 2400.670 ;
        RECT 775.730 2399.490 776.910 2400.670 ;
        RECT 774.130 2221.090 775.310 2222.270 ;
        RECT 775.730 2221.090 776.910 2222.270 ;
        RECT 774.130 2219.490 775.310 2220.670 ;
        RECT 775.730 2219.490 776.910 2220.670 ;
        RECT 774.130 2041.090 775.310 2042.270 ;
        RECT 775.730 2041.090 776.910 2042.270 ;
        RECT 774.130 2039.490 775.310 2040.670 ;
        RECT 775.730 2039.490 776.910 2040.670 ;
        RECT 774.130 1861.090 775.310 1862.270 ;
        RECT 775.730 1861.090 776.910 1862.270 ;
        RECT 774.130 1859.490 775.310 1860.670 ;
        RECT 775.730 1859.490 776.910 1860.670 ;
        RECT 774.130 1681.090 775.310 1682.270 ;
        RECT 775.730 1681.090 776.910 1682.270 ;
        RECT 774.130 1679.490 775.310 1680.670 ;
        RECT 775.730 1679.490 776.910 1680.670 ;
        RECT 774.130 1501.090 775.310 1502.270 ;
        RECT 775.730 1501.090 776.910 1502.270 ;
        RECT 774.130 1499.490 775.310 1500.670 ;
        RECT 775.730 1499.490 776.910 1500.670 ;
        RECT 774.130 1321.090 775.310 1322.270 ;
        RECT 775.730 1321.090 776.910 1322.270 ;
        RECT 774.130 1319.490 775.310 1320.670 ;
        RECT 775.730 1319.490 776.910 1320.670 ;
        RECT 774.130 1141.090 775.310 1142.270 ;
        RECT 775.730 1141.090 776.910 1142.270 ;
        RECT 774.130 1139.490 775.310 1140.670 ;
        RECT 775.730 1139.490 776.910 1140.670 ;
        RECT 774.130 961.090 775.310 962.270 ;
        RECT 775.730 961.090 776.910 962.270 ;
        RECT 774.130 959.490 775.310 960.670 ;
        RECT 775.730 959.490 776.910 960.670 ;
        RECT 234.130 781.090 235.310 782.270 ;
        RECT 235.730 781.090 236.910 782.270 ;
        RECT 234.130 779.490 235.310 780.670 ;
        RECT 235.730 779.490 236.910 780.670 ;
        RECT 234.130 601.090 235.310 602.270 ;
        RECT 235.730 601.090 236.910 602.270 ;
        RECT 234.130 599.490 235.310 600.670 ;
        RECT 235.730 599.490 236.910 600.670 ;
        RECT 774.130 781.090 775.310 782.270 ;
        RECT 775.730 781.090 776.910 782.270 ;
        RECT 774.130 779.490 775.310 780.670 ;
        RECT 775.730 779.490 776.910 780.670 ;
        RECT 774.130 601.090 775.310 602.270 ;
        RECT 775.730 601.090 776.910 602.270 ;
        RECT 774.130 599.490 775.310 600.670 ;
        RECT 775.730 599.490 776.910 600.670 ;
        RECT 234.130 421.090 235.310 422.270 ;
        RECT 235.730 421.090 236.910 422.270 ;
        RECT 234.130 419.490 235.310 420.670 ;
        RECT 235.730 419.490 236.910 420.670 ;
        RECT 234.130 241.090 235.310 242.270 ;
        RECT 235.730 241.090 236.910 242.270 ;
        RECT 234.130 239.490 235.310 240.670 ;
        RECT 235.730 239.490 236.910 240.670 ;
        RECT 234.130 61.090 235.310 62.270 ;
        RECT 235.730 61.090 236.910 62.270 ;
        RECT 234.130 59.490 235.310 60.670 ;
        RECT 235.730 59.490 236.910 60.670 ;
        RECT 234.130 -12.510 235.310 -11.330 ;
        RECT 235.730 -12.510 236.910 -11.330 ;
        RECT 234.130 -14.110 235.310 -12.930 ;
        RECT 235.730 -14.110 236.910 -12.930 ;
        RECT 414.130 421.090 415.310 422.270 ;
        RECT 415.730 421.090 416.910 422.270 ;
        RECT 414.130 419.490 415.310 420.670 ;
        RECT 415.730 419.490 416.910 420.670 ;
        RECT 414.130 241.090 415.310 242.270 ;
        RECT 415.730 241.090 416.910 242.270 ;
        RECT 414.130 239.490 415.310 240.670 ;
        RECT 415.730 239.490 416.910 240.670 ;
        RECT 414.130 61.090 415.310 62.270 ;
        RECT 415.730 61.090 416.910 62.270 ;
        RECT 414.130 59.490 415.310 60.670 ;
        RECT 415.730 59.490 416.910 60.670 ;
        RECT 414.130 -12.510 415.310 -11.330 ;
        RECT 415.730 -12.510 416.910 -11.330 ;
        RECT 414.130 -14.110 415.310 -12.930 ;
        RECT 415.730 -14.110 416.910 -12.930 ;
        RECT 594.130 421.090 595.310 422.270 ;
        RECT 595.730 421.090 596.910 422.270 ;
        RECT 594.130 419.490 595.310 420.670 ;
        RECT 595.730 419.490 596.910 420.670 ;
        RECT 594.130 241.090 595.310 242.270 ;
        RECT 595.730 241.090 596.910 242.270 ;
        RECT 594.130 239.490 595.310 240.670 ;
        RECT 595.730 239.490 596.910 240.670 ;
        RECT 594.130 61.090 595.310 62.270 ;
        RECT 595.730 61.090 596.910 62.270 ;
        RECT 594.130 59.490 595.310 60.670 ;
        RECT 595.730 59.490 596.910 60.670 ;
        RECT 594.130 -12.510 595.310 -11.330 ;
        RECT 595.730 -12.510 596.910 -11.330 ;
        RECT 594.130 -14.110 595.310 -12.930 ;
        RECT 595.730 -14.110 596.910 -12.930 ;
        RECT 774.130 421.090 775.310 422.270 ;
        RECT 775.730 421.090 776.910 422.270 ;
        RECT 774.130 419.490 775.310 420.670 ;
        RECT 775.730 419.490 776.910 420.670 ;
        RECT 774.130 241.090 775.310 242.270 ;
        RECT 775.730 241.090 776.910 242.270 ;
        RECT 774.130 239.490 775.310 240.670 ;
        RECT 775.730 239.490 776.910 240.670 ;
        RECT 774.130 61.090 775.310 62.270 ;
        RECT 775.730 61.090 776.910 62.270 ;
        RECT 774.130 59.490 775.310 60.670 ;
        RECT 775.730 59.490 776.910 60.670 ;
        RECT 774.130 -12.510 775.310 -11.330 ;
        RECT 775.730 -12.510 776.910 -11.330 ;
        RECT 774.130 -14.110 775.310 -12.930 ;
        RECT 775.730 -14.110 776.910 -12.930 ;
        RECT 954.130 3532.610 955.310 3533.790 ;
        RECT 955.730 3532.610 956.910 3533.790 ;
        RECT 954.130 3531.010 955.310 3532.190 ;
        RECT 955.730 3531.010 956.910 3532.190 ;
        RECT 954.130 3481.090 955.310 3482.270 ;
        RECT 955.730 3481.090 956.910 3482.270 ;
        RECT 954.130 3479.490 955.310 3480.670 ;
        RECT 955.730 3479.490 956.910 3480.670 ;
        RECT 954.130 3301.090 955.310 3302.270 ;
        RECT 955.730 3301.090 956.910 3302.270 ;
        RECT 954.130 3299.490 955.310 3300.670 ;
        RECT 955.730 3299.490 956.910 3300.670 ;
        RECT 954.130 3121.090 955.310 3122.270 ;
        RECT 955.730 3121.090 956.910 3122.270 ;
        RECT 954.130 3119.490 955.310 3120.670 ;
        RECT 955.730 3119.490 956.910 3120.670 ;
        RECT 954.130 2941.090 955.310 2942.270 ;
        RECT 955.730 2941.090 956.910 2942.270 ;
        RECT 954.130 2939.490 955.310 2940.670 ;
        RECT 955.730 2939.490 956.910 2940.670 ;
        RECT 954.130 2761.090 955.310 2762.270 ;
        RECT 955.730 2761.090 956.910 2762.270 ;
        RECT 954.130 2759.490 955.310 2760.670 ;
        RECT 955.730 2759.490 956.910 2760.670 ;
        RECT 954.130 2581.090 955.310 2582.270 ;
        RECT 955.730 2581.090 956.910 2582.270 ;
        RECT 954.130 2579.490 955.310 2580.670 ;
        RECT 955.730 2579.490 956.910 2580.670 ;
        RECT 954.130 2401.090 955.310 2402.270 ;
        RECT 955.730 2401.090 956.910 2402.270 ;
        RECT 954.130 2399.490 955.310 2400.670 ;
        RECT 955.730 2399.490 956.910 2400.670 ;
        RECT 954.130 2221.090 955.310 2222.270 ;
        RECT 955.730 2221.090 956.910 2222.270 ;
        RECT 954.130 2219.490 955.310 2220.670 ;
        RECT 955.730 2219.490 956.910 2220.670 ;
        RECT 954.130 2041.090 955.310 2042.270 ;
        RECT 955.730 2041.090 956.910 2042.270 ;
        RECT 954.130 2039.490 955.310 2040.670 ;
        RECT 955.730 2039.490 956.910 2040.670 ;
        RECT 954.130 1861.090 955.310 1862.270 ;
        RECT 955.730 1861.090 956.910 1862.270 ;
        RECT 954.130 1859.490 955.310 1860.670 ;
        RECT 955.730 1859.490 956.910 1860.670 ;
        RECT 954.130 1681.090 955.310 1682.270 ;
        RECT 955.730 1681.090 956.910 1682.270 ;
        RECT 954.130 1679.490 955.310 1680.670 ;
        RECT 955.730 1679.490 956.910 1680.670 ;
        RECT 954.130 1501.090 955.310 1502.270 ;
        RECT 955.730 1501.090 956.910 1502.270 ;
        RECT 954.130 1499.490 955.310 1500.670 ;
        RECT 955.730 1499.490 956.910 1500.670 ;
        RECT 954.130 1321.090 955.310 1322.270 ;
        RECT 955.730 1321.090 956.910 1322.270 ;
        RECT 954.130 1319.490 955.310 1320.670 ;
        RECT 955.730 1319.490 956.910 1320.670 ;
        RECT 954.130 1141.090 955.310 1142.270 ;
        RECT 955.730 1141.090 956.910 1142.270 ;
        RECT 954.130 1139.490 955.310 1140.670 ;
        RECT 955.730 1139.490 956.910 1140.670 ;
        RECT 954.130 961.090 955.310 962.270 ;
        RECT 955.730 961.090 956.910 962.270 ;
        RECT 954.130 959.490 955.310 960.670 ;
        RECT 955.730 959.490 956.910 960.670 ;
        RECT 954.130 781.090 955.310 782.270 ;
        RECT 955.730 781.090 956.910 782.270 ;
        RECT 954.130 779.490 955.310 780.670 ;
        RECT 955.730 779.490 956.910 780.670 ;
        RECT 954.130 601.090 955.310 602.270 ;
        RECT 955.730 601.090 956.910 602.270 ;
        RECT 954.130 599.490 955.310 600.670 ;
        RECT 955.730 599.490 956.910 600.670 ;
        RECT 954.130 421.090 955.310 422.270 ;
        RECT 955.730 421.090 956.910 422.270 ;
        RECT 954.130 419.490 955.310 420.670 ;
        RECT 955.730 419.490 956.910 420.670 ;
        RECT 954.130 241.090 955.310 242.270 ;
        RECT 955.730 241.090 956.910 242.270 ;
        RECT 954.130 239.490 955.310 240.670 ;
        RECT 955.730 239.490 956.910 240.670 ;
        RECT 954.130 61.090 955.310 62.270 ;
        RECT 955.730 61.090 956.910 62.270 ;
        RECT 954.130 59.490 955.310 60.670 ;
        RECT 955.730 59.490 956.910 60.670 ;
        RECT 954.130 -12.510 955.310 -11.330 ;
        RECT 955.730 -12.510 956.910 -11.330 ;
        RECT 954.130 -14.110 955.310 -12.930 ;
        RECT 955.730 -14.110 956.910 -12.930 ;
        RECT 1134.130 3532.610 1135.310 3533.790 ;
        RECT 1135.730 3532.610 1136.910 3533.790 ;
        RECT 1134.130 3531.010 1135.310 3532.190 ;
        RECT 1135.730 3531.010 1136.910 3532.190 ;
        RECT 1134.130 3481.090 1135.310 3482.270 ;
        RECT 1135.730 3481.090 1136.910 3482.270 ;
        RECT 1134.130 3479.490 1135.310 3480.670 ;
        RECT 1135.730 3479.490 1136.910 3480.670 ;
        RECT 1134.130 3301.090 1135.310 3302.270 ;
        RECT 1135.730 3301.090 1136.910 3302.270 ;
        RECT 1134.130 3299.490 1135.310 3300.670 ;
        RECT 1135.730 3299.490 1136.910 3300.670 ;
        RECT 1134.130 3121.090 1135.310 3122.270 ;
        RECT 1135.730 3121.090 1136.910 3122.270 ;
        RECT 1134.130 3119.490 1135.310 3120.670 ;
        RECT 1135.730 3119.490 1136.910 3120.670 ;
        RECT 1134.130 2941.090 1135.310 2942.270 ;
        RECT 1135.730 2941.090 1136.910 2942.270 ;
        RECT 1134.130 2939.490 1135.310 2940.670 ;
        RECT 1135.730 2939.490 1136.910 2940.670 ;
        RECT 1134.130 2761.090 1135.310 2762.270 ;
        RECT 1135.730 2761.090 1136.910 2762.270 ;
        RECT 1134.130 2759.490 1135.310 2760.670 ;
        RECT 1135.730 2759.490 1136.910 2760.670 ;
        RECT 1134.130 2581.090 1135.310 2582.270 ;
        RECT 1135.730 2581.090 1136.910 2582.270 ;
        RECT 1134.130 2579.490 1135.310 2580.670 ;
        RECT 1135.730 2579.490 1136.910 2580.670 ;
        RECT 1134.130 2401.090 1135.310 2402.270 ;
        RECT 1135.730 2401.090 1136.910 2402.270 ;
        RECT 1134.130 2399.490 1135.310 2400.670 ;
        RECT 1135.730 2399.490 1136.910 2400.670 ;
        RECT 1134.130 2221.090 1135.310 2222.270 ;
        RECT 1135.730 2221.090 1136.910 2222.270 ;
        RECT 1134.130 2219.490 1135.310 2220.670 ;
        RECT 1135.730 2219.490 1136.910 2220.670 ;
        RECT 1134.130 2041.090 1135.310 2042.270 ;
        RECT 1135.730 2041.090 1136.910 2042.270 ;
        RECT 1134.130 2039.490 1135.310 2040.670 ;
        RECT 1135.730 2039.490 1136.910 2040.670 ;
        RECT 1134.130 1861.090 1135.310 1862.270 ;
        RECT 1135.730 1861.090 1136.910 1862.270 ;
        RECT 1134.130 1859.490 1135.310 1860.670 ;
        RECT 1135.730 1859.490 1136.910 1860.670 ;
        RECT 1134.130 1681.090 1135.310 1682.270 ;
        RECT 1135.730 1681.090 1136.910 1682.270 ;
        RECT 1134.130 1679.490 1135.310 1680.670 ;
        RECT 1135.730 1679.490 1136.910 1680.670 ;
        RECT 1134.130 1501.090 1135.310 1502.270 ;
        RECT 1135.730 1501.090 1136.910 1502.270 ;
        RECT 1134.130 1499.490 1135.310 1500.670 ;
        RECT 1135.730 1499.490 1136.910 1500.670 ;
        RECT 1134.130 1321.090 1135.310 1322.270 ;
        RECT 1135.730 1321.090 1136.910 1322.270 ;
        RECT 1134.130 1319.490 1135.310 1320.670 ;
        RECT 1135.730 1319.490 1136.910 1320.670 ;
        RECT 1134.130 1141.090 1135.310 1142.270 ;
        RECT 1135.730 1141.090 1136.910 1142.270 ;
        RECT 1134.130 1139.490 1135.310 1140.670 ;
        RECT 1135.730 1139.490 1136.910 1140.670 ;
        RECT 1134.130 961.090 1135.310 962.270 ;
        RECT 1135.730 961.090 1136.910 962.270 ;
        RECT 1134.130 959.490 1135.310 960.670 ;
        RECT 1135.730 959.490 1136.910 960.670 ;
        RECT 1134.130 781.090 1135.310 782.270 ;
        RECT 1135.730 781.090 1136.910 782.270 ;
        RECT 1134.130 779.490 1135.310 780.670 ;
        RECT 1135.730 779.490 1136.910 780.670 ;
        RECT 1134.130 601.090 1135.310 602.270 ;
        RECT 1135.730 601.090 1136.910 602.270 ;
        RECT 1134.130 599.490 1135.310 600.670 ;
        RECT 1135.730 599.490 1136.910 600.670 ;
        RECT 1134.130 421.090 1135.310 422.270 ;
        RECT 1135.730 421.090 1136.910 422.270 ;
        RECT 1134.130 419.490 1135.310 420.670 ;
        RECT 1135.730 419.490 1136.910 420.670 ;
        RECT 1134.130 241.090 1135.310 242.270 ;
        RECT 1135.730 241.090 1136.910 242.270 ;
        RECT 1134.130 239.490 1135.310 240.670 ;
        RECT 1135.730 239.490 1136.910 240.670 ;
        RECT 1134.130 61.090 1135.310 62.270 ;
        RECT 1135.730 61.090 1136.910 62.270 ;
        RECT 1134.130 59.490 1135.310 60.670 ;
        RECT 1135.730 59.490 1136.910 60.670 ;
        RECT 1134.130 -12.510 1135.310 -11.330 ;
        RECT 1135.730 -12.510 1136.910 -11.330 ;
        RECT 1134.130 -14.110 1135.310 -12.930 ;
        RECT 1135.730 -14.110 1136.910 -12.930 ;
        RECT 1314.130 3532.610 1315.310 3533.790 ;
        RECT 1315.730 3532.610 1316.910 3533.790 ;
        RECT 1314.130 3531.010 1315.310 3532.190 ;
        RECT 1315.730 3531.010 1316.910 3532.190 ;
        RECT 1314.130 3481.090 1315.310 3482.270 ;
        RECT 1315.730 3481.090 1316.910 3482.270 ;
        RECT 1314.130 3479.490 1315.310 3480.670 ;
        RECT 1315.730 3479.490 1316.910 3480.670 ;
        RECT 1314.130 3301.090 1315.310 3302.270 ;
        RECT 1315.730 3301.090 1316.910 3302.270 ;
        RECT 1314.130 3299.490 1315.310 3300.670 ;
        RECT 1315.730 3299.490 1316.910 3300.670 ;
        RECT 1314.130 3121.090 1315.310 3122.270 ;
        RECT 1315.730 3121.090 1316.910 3122.270 ;
        RECT 1314.130 3119.490 1315.310 3120.670 ;
        RECT 1315.730 3119.490 1316.910 3120.670 ;
        RECT 1314.130 2941.090 1315.310 2942.270 ;
        RECT 1315.730 2941.090 1316.910 2942.270 ;
        RECT 1314.130 2939.490 1315.310 2940.670 ;
        RECT 1315.730 2939.490 1316.910 2940.670 ;
        RECT 1314.130 2761.090 1315.310 2762.270 ;
        RECT 1315.730 2761.090 1316.910 2762.270 ;
        RECT 1314.130 2759.490 1315.310 2760.670 ;
        RECT 1315.730 2759.490 1316.910 2760.670 ;
        RECT 1314.130 2581.090 1315.310 2582.270 ;
        RECT 1315.730 2581.090 1316.910 2582.270 ;
        RECT 1314.130 2579.490 1315.310 2580.670 ;
        RECT 1315.730 2579.490 1316.910 2580.670 ;
        RECT 1314.130 2401.090 1315.310 2402.270 ;
        RECT 1315.730 2401.090 1316.910 2402.270 ;
        RECT 1314.130 2399.490 1315.310 2400.670 ;
        RECT 1315.730 2399.490 1316.910 2400.670 ;
        RECT 1314.130 2221.090 1315.310 2222.270 ;
        RECT 1315.730 2221.090 1316.910 2222.270 ;
        RECT 1314.130 2219.490 1315.310 2220.670 ;
        RECT 1315.730 2219.490 1316.910 2220.670 ;
        RECT 1314.130 2041.090 1315.310 2042.270 ;
        RECT 1315.730 2041.090 1316.910 2042.270 ;
        RECT 1314.130 2039.490 1315.310 2040.670 ;
        RECT 1315.730 2039.490 1316.910 2040.670 ;
        RECT 1314.130 1861.090 1315.310 1862.270 ;
        RECT 1315.730 1861.090 1316.910 1862.270 ;
        RECT 1314.130 1859.490 1315.310 1860.670 ;
        RECT 1315.730 1859.490 1316.910 1860.670 ;
        RECT 1314.130 1681.090 1315.310 1682.270 ;
        RECT 1315.730 1681.090 1316.910 1682.270 ;
        RECT 1314.130 1679.490 1315.310 1680.670 ;
        RECT 1315.730 1679.490 1316.910 1680.670 ;
        RECT 1314.130 1501.090 1315.310 1502.270 ;
        RECT 1315.730 1501.090 1316.910 1502.270 ;
        RECT 1314.130 1499.490 1315.310 1500.670 ;
        RECT 1315.730 1499.490 1316.910 1500.670 ;
        RECT 1314.130 1321.090 1315.310 1322.270 ;
        RECT 1315.730 1321.090 1316.910 1322.270 ;
        RECT 1314.130 1319.490 1315.310 1320.670 ;
        RECT 1315.730 1319.490 1316.910 1320.670 ;
        RECT 1314.130 1141.090 1315.310 1142.270 ;
        RECT 1315.730 1141.090 1316.910 1142.270 ;
        RECT 1314.130 1139.490 1315.310 1140.670 ;
        RECT 1315.730 1139.490 1316.910 1140.670 ;
        RECT 1314.130 961.090 1315.310 962.270 ;
        RECT 1315.730 961.090 1316.910 962.270 ;
        RECT 1314.130 959.490 1315.310 960.670 ;
        RECT 1315.730 959.490 1316.910 960.670 ;
        RECT 1314.130 781.090 1315.310 782.270 ;
        RECT 1315.730 781.090 1316.910 782.270 ;
        RECT 1314.130 779.490 1315.310 780.670 ;
        RECT 1315.730 779.490 1316.910 780.670 ;
        RECT 1314.130 601.090 1315.310 602.270 ;
        RECT 1315.730 601.090 1316.910 602.270 ;
        RECT 1314.130 599.490 1315.310 600.670 ;
        RECT 1315.730 599.490 1316.910 600.670 ;
        RECT 1314.130 421.090 1315.310 422.270 ;
        RECT 1315.730 421.090 1316.910 422.270 ;
        RECT 1314.130 419.490 1315.310 420.670 ;
        RECT 1315.730 419.490 1316.910 420.670 ;
        RECT 1314.130 241.090 1315.310 242.270 ;
        RECT 1315.730 241.090 1316.910 242.270 ;
        RECT 1314.130 239.490 1315.310 240.670 ;
        RECT 1315.730 239.490 1316.910 240.670 ;
        RECT 1314.130 61.090 1315.310 62.270 ;
        RECT 1315.730 61.090 1316.910 62.270 ;
        RECT 1314.130 59.490 1315.310 60.670 ;
        RECT 1315.730 59.490 1316.910 60.670 ;
        RECT 1314.130 -12.510 1315.310 -11.330 ;
        RECT 1315.730 -12.510 1316.910 -11.330 ;
        RECT 1314.130 -14.110 1315.310 -12.930 ;
        RECT 1315.730 -14.110 1316.910 -12.930 ;
        RECT 1494.130 3532.610 1495.310 3533.790 ;
        RECT 1495.730 3532.610 1496.910 3533.790 ;
        RECT 1494.130 3531.010 1495.310 3532.190 ;
        RECT 1495.730 3531.010 1496.910 3532.190 ;
        RECT 1494.130 3481.090 1495.310 3482.270 ;
        RECT 1495.730 3481.090 1496.910 3482.270 ;
        RECT 1494.130 3479.490 1495.310 3480.670 ;
        RECT 1495.730 3479.490 1496.910 3480.670 ;
        RECT 1494.130 3301.090 1495.310 3302.270 ;
        RECT 1495.730 3301.090 1496.910 3302.270 ;
        RECT 1494.130 3299.490 1495.310 3300.670 ;
        RECT 1495.730 3299.490 1496.910 3300.670 ;
        RECT 1494.130 3121.090 1495.310 3122.270 ;
        RECT 1495.730 3121.090 1496.910 3122.270 ;
        RECT 1494.130 3119.490 1495.310 3120.670 ;
        RECT 1495.730 3119.490 1496.910 3120.670 ;
        RECT 1494.130 2941.090 1495.310 2942.270 ;
        RECT 1495.730 2941.090 1496.910 2942.270 ;
        RECT 1494.130 2939.490 1495.310 2940.670 ;
        RECT 1495.730 2939.490 1496.910 2940.670 ;
        RECT 1494.130 2761.090 1495.310 2762.270 ;
        RECT 1495.730 2761.090 1496.910 2762.270 ;
        RECT 1494.130 2759.490 1495.310 2760.670 ;
        RECT 1495.730 2759.490 1496.910 2760.670 ;
        RECT 1494.130 2581.090 1495.310 2582.270 ;
        RECT 1495.730 2581.090 1496.910 2582.270 ;
        RECT 1494.130 2579.490 1495.310 2580.670 ;
        RECT 1495.730 2579.490 1496.910 2580.670 ;
        RECT 1494.130 2401.090 1495.310 2402.270 ;
        RECT 1495.730 2401.090 1496.910 2402.270 ;
        RECT 1494.130 2399.490 1495.310 2400.670 ;
        RECT 1495.730 2399.490 1496.910 2400.670 ;
        RECT 1494.130 2221.090 1495.310 2222.270 ;
        RECT 1495.730 2221.090 1496.910 2222.270 ;
        RECT 1494.130 2219.490 1495.310 2220.670 ;
        RECT 1495.730 2219.490 1496.910 2220.670 ;
        RECT 1494.130 2041.090 1495.310 2042.270 ;
        RECT 1495.730 2041.090 1496.910 2042.270 ;
        RECT 1494.130 2039.490 1495.310 2040.670 ;
        RECT 1495.730 2039.490 1496.910 2040.670 ;
        RECT 1494.130 1861.090 1495.310 1862.270 ;
        RECT 1495.730 1861.090 1496.910 1862.270 ;
        RECT 1494.130 1859.490 1495.310 1860.670 ;
        RECT 1495.730 1859.490 1496.910 1860.670 ;
        RECT 1494.130 1681.090 1495.310 1682.270 ;
        RECT 1495.730 1681.090 1496.910 1682.270 ;
        RECT 1494.130 1679.490 1495.310 1680.670 ;
        RECT 1495.730 1679.490 1496.910 1680.670 ;
        RECT 1494.130 1501.090 1495.310 1502.270 ;
        RECT 1495.730 1501.090 1496.910 1502.270 ;
        RECT 1494.130 1499.490 1495.310 1500.670 ;
        RECT 1495.730 1499.490 1496.910 1500.670 ;
        RECT 1494.130 1321.090 1495.310 1322.270 ;
        RECT 1495.730 1321.090 1496.910 1322.270 ;
        RECT 1494.130 1319.490 1495.310 1320.670 ;
        RECT 1495.730 1319.490 1496.910 1320.670 ;
        RECT 1494.130 1141.090 1495.310 1142.270 ;
        RECT 1495.730 1141.090 1496.910 1142.270 ;
        RECT 1494.130 1139.490 1495.310 1140.670 ;
        RECT 1495.730 1139.490 1496.910 1140.670 ;
        RECT 1494.130 961.090 1495.310 962.270 ;
        RECT 1495.730 961.090 1496.910 962.270 ;
        RECT 1494.130 959.490 1495.310 960.670 ;
        RECT 1495.730 959.490 1496.910 960.670 ;
        RECT 1494.130 781.090 1495.310 782.270 ;
        RECT 1495.730 781.090 1496.910 782.270 ;
        RECT 1494.130 779.490 1495.310 780.670 ;
        RECT 1495.730 779.490 1496.910 780.670 ;
        RECT 1494.130 601.090 1495.310 602.270 ;
        RECT 1495.730 601.090 1496.910 602.270 ;
        RECT 1494.130 599.490 1495.310 600.670 ;
        RECT 1495.730 599.490 1496.910 600.670 ;
        RECT 1494.130 421.090 1495.310 422.270 ;
        RECT 1495.730 421.090 1496.910 422.270 ;
        RECT 1494.130 419.490 1495.310 420.670 ;
        RECT 1495.730 419.490 1496.910 420.670 ;
        RECT 1494.130 241.090 1495.310 242.270 ;
        RECT 1495.730 241.090 1496.910 242.270 ;
        RECT 1494.130 239.490 1495.310 240.670 ;
        RECT 1495.730 239.490 1496.910 240.670 ;
        RECT 1494.130 61.090 1495.310 62.270 ;
        RECT 1495.730 61.090 1496.910 62.270 ;
        RECT 1494.130 59.490 1495.310 60.670 ;
        RECT 1495.730 59.490 1496.910 60.670 ;
        RECT 1494.130 -12.510 1495.310 -11.330 ;
        RECT 1495.730 -12.510 1496.910 -11.330 ;
        RECT 1494.130 -14.110 1495.310 -12.930 ;
        RECT 1495.730 -14.110 1496.910 -12.930 ;
        RECT 1674.130 3532.610 1675.310 3533.790 ;
        RECT 1675.730 3532.610 1676.910 3533.790 ;
        RECT 1674.130 3531.010 1675.310 3532.190 ;
        RECT 1675.730 3531.010 1676.910 3532.190 ;
        RECT 1674.130 3481.090 1675.310 3482.270 ;
        RECT 1675.730 3481.090 1676.910 3482.270 ;
        RECT 1674.130 3479.490 1675.310 3480.670 ;
        RECT 1675.730 3479.490 1676.910 3480.670 ;
        RECT 1674.130 3301.090 1675.310 3302.270 ;
        RECT 1675.730 3301.090 1676.910 3302.270 ;
        RECT 1674.130 3299.490 1675.310 3300.670 ;
        RECT 1675.730 3299.490 1676.910 3300.670 ;
        RECT 1674.130 3121.090 1675.310 3122.270 ;
        RECT 1675.730 3121.090 1676.910 3122.270 ;
        RECT 1674.130 3119.490 1675.310 3120.670 ;
        RECT 1675.730 3119.490 1676.910 3120.670 ;
        RECT 1674.130 2941.090 1675.310 2942.270 ;
        RECT 1675.730 2941.090 1676.910 2942.270 ;
        RECT 1674.130 2939.490 1675.310 2940.670 ;
        RECT 1675.730 2939.490 1676.910 2940.670 ;
        RECT 1674.130 2761.090 1675.310 2762.270 ;
        RECT 1675.730 2761.090 1676.910 2762.270 ;
        RECT 1674.130 2759.490 1675.310 2760.670 ;
        RECT 1675.730 2759.490 1676.910 2760.670 ;
        RECT 1674.130 2581.090 1675.310 2582.270 ;
        RECT 1675.730 2581.090 1676.910 2582.270 ;
        RECT 1674.130 2579.490 1675.310 2580.670 ;
        RECT 1675.730 2579.490 1676.910 2580.670 ;
        RECT 1674.130 2401.090 1675.310 2402.270 ;
        RECT 1675.730 2401.090 1676.910 2402.270 ;
        RECT 1674.130 2399.490 1675.310 2400.670 ;
        RECT 1675.730 2399.490 1676.910 2400.670 ;
        RECT 1674.130 2221.090 1675.310 2222.270 ;
        RECT 1675.730 2221.090 1676.910 2222.270 ;
        RECT 1674.130 2219.490 1675.310 2220.670 ;
        RECT 1675.730 2219.490 1676.910 2220.670 ;
        RECT 1674.130 2041.090 1675.310 2042.270 ;
        RECT 1675.730 2041.090 1676.910 2042.270 ;
        RECT 1674.130 2039.490 1675.310 2040.670 ;
        RECT 1675.730 2039.490 1676.910 2040.670 ;
        RECT 1674.130 1861.090 1675.310 1862.270 ;
        RECT 1675.730 1861.090 1676.910 1862.270 ;
        RECT 1674.130 1859.490 1675.310 1860.670 ;
        RECT 1675.730 1859.490 1676.910 1860.670 ;
        RECT 1674.130 1681.090 1675.310 1682.270 ;
        RECT 1675.730 1681.090 1676.910 1682.270 ;
        RECT 1674.130 1679.490 1675.310 1680.670 ;
        RECT 1675.730 1679.490 1676.910 1680.670 ;
        RECT 1674.130 1501.090 1675.310 1502.270 ;
        RECT 1675.730 1501.090 1676.910 1502.270 ;
        RECT 1674.130 1499.490 1675.310 1500.670 ;
        RECT 1675.730 1499.490 1676.910 1500.670 ;
        RECT 1674.130 1321.090 1675.310 1322.270 ;
        RECT 1675.730 1321.090 1676.910 1322.270 ;
        RECT 1674.130 1319.490 1675.310 1320.670 ;
        RECT 1675.730 1319.490 1676.910 1320.670 ;
        RECT 1674.130 1141.090 1675.310 1142.270 ;
        RECT 1675.730 1141.090 1676.910 1142.270 ;
        RECT 1674.130 1139.490 1675.310 1140.670 ;
        RECT 1675.730 1139.490 1676.910 1140.670 ;
        RECT 1674.130 961.090 1675.310 962.270 ;
        RECT 1675.730 961.090 1676.910 962.270 ;
        RECT 1674.130 959.490 1675.310 960.670 ;
        RECT 1675.730 959.490 1676.910 960.670 ;
        RECT 1674.130 781.090 1675.310 782.270 ;
        RECT 1675.730 781.090 1676.910 782.270 ;
        RECT 1674.130 779.490 1675.310 780.670 ;
        RECT 1675.730 779.490 1676.910 780.670 ;
        RECT 1674.130 601.090 1675.310 602.270 ;
        RECT 1675.730 601.090 1676.910 602.270 ;
        RECT 1674.130 599.490 1675.310 600.670 ;
        RECT 1675.730 599.490 1676.910 600.670 ;
        RECT 1674.130 421.090 1675.310 422.270 ;
        RECT 1675.730 421.090 1676.910 422.270 ;
        RECT 1674.130 419.490 1675.310 420.670 ;
        RECT 1675.730 419.490 1676.910 420.670 ;
        RECT 1674.130 241.090 1675.310 242.270 ;
        RECT 1675.730 241.090 1676.910 242.270 ;
        RECT 1674.130 239.490 1675.310 240.670 ;
        RECT 1675.730 239.490 1676.910 240.670 ;
        RECT 1674.130 61.090 1675.310 62.270 ;
        RECT 1675.730 61.090 1676.910 62.270 ;
        RECT 1674.130 59.490 1675.310 60.670 ;
        RECT 1675.730 59.490 1676.910 60.670 ;
        RECT 1674.130 -12.510 1675.310 -11.330 ;
        RECT 1675.730 -12.510 1676.910 -11.330 ;
        RECT 1674.130 -14.110 1675.310 -12.930 ;
        RECT 1675.730 -14.110 1676.910 -12.930 ;
        RECT 1854.130 3532.610 1855.310 3533.790 ;
        RECT 1855.730 3532.610 1856.910 3533.790 ;
        RECT 1854.130 3531.010 1855.310 3532.190 ;
        RECT 1855.730 3531.010 1856.910 3532.190 ;
        RECT 1854.130 3481.090 1855.310 3482.270 ;
        RECT 1855.730 3481.090 1856.910 3482.270 ;
        RECT 1854.130 3479.490 1855.310 3480.670 ;
        RECT 1855.730 3479.490 1856.910 3480.670 ;
        RECT 1854.130 3301.090 1855.310 3302.270 ;
        RECT 1855.730 3301.090 1856.910 3302.270 ;
        RECT 1854.130 3299.490 1855.310 3300.670 ;
        RECT 1855.730 3299.490 1856.910 3300.670 ;
        RECT 1854.130 3121.090 1855.310 3122.270 ;
        RECT 1855.730 3121.090 1856.910 3122.270 ;
        RECT 1854.130 3119.490 1855.310 3120.670 ;
        RECT 1855.730 3119.490 1856.910 3120.670 ;
        RECT 1854.130 2941.090 1855.310 2942.270 ;
        RECT 1855.730 2941.090 1856.910 2942.270 ;
        RECT 1854.130 2939.490 1855.310 2940.670 ;
        RECT 1855.730 2939.490 1856.910 2940.670 ;
        RECT 1854.130 2761.090 1855.310 2762.270 ;
        RECT 1855.730 2761.090 1856.910 2762.270 ;
        RECT 1854.130 2759.490 1855.310 2760.670 ;
        RECT 1855.730 2759.490 1856.910 2760.670 ;
        RECT 1854.130 2581.090 1855.310 2582.270 ;
        RECT 1855.730 2581.090 1856.910 2582.270 ;
        RECT 1854.130 2579.490 1855.310 2580.670 ;
        RECT 1855.730 2579.490 1856.910 2580.670 ;
        RECT 1854.130 2401.090 1855.310 2402.270 ;
        RECT 1855.730 2401.090 1856.910 2402.270 ;
        RECT 1854.130 2399.490 1855.310 2400.670 ;
        RECT 1855.730 2399.490 1856.910 2400.670 ;
        RECT 1854.130 2221.090 1855.310 2222.270 ;
        RECT 1855.730 2221.090 1856.910 2222.270 ;
        RECT 1854.130 2219.490 1855.310 2220.670 ;
        RECT 1855.730 2219.490 1856.910 2220.670 ;
        RECT 1854.130 2041.090 1855.310 2042.270 ;
        RECT 1855.730 2041.090 1856.910 2042.270 ;
        RECT 1854.130 2039.490 1855.310 2040.670 ;
        RECT 1855.730 2039.490 1856.910 2040.670 ;
        RECT 1854.130 1861.090 1855.310 1862.270 ;
        RECT 1855.730 1861.090 1856.910 1862.270 ;
        RECT 1854.130 1859.490 1855.310 1860.670 ;
        RECT 1855.730 1859.490 1856.910 1860.670 ;
        RECT 1854.130 1681.090 1855.310 1682.270 ;
        RECT 1855.730 1681.090 1856.910 1682.270 ;
        RECT 1854.130 1679.490 1855.310 1680.670 ;
        RECT 1855.730 1679.490 1856.910 1680.670 ;
        RECT 1854.130 1501.090 1855.310 1502.270 ;
        RECT 1855.730 1501.090 1856.910 1502.270 ;
        RECT 1854.130 1499.490 1855.310 1500.670 ;
        RECT 1855.730 1499.490 1856.910 1500.670 ;
        RECT 1854.130 1321.090 1855.310 1322.270 ;
        RECT 1855.730 1321.090 1856.910 1322.270 ;
        RECT 1854.130 1319.490 1855.310 1320.670 ;
        RECT 1855.730 1319.490 1856.910 1320.670 ;
        RECT 1854.130 1141.090 1855.310 1142.270 ;
        RECT 1855.730 1141.090 1856.910 1142.270 ;
        RECT 1854.130 1139.490 1855.310 1140.670 ;
        RECT 1855.730 1139.490 1856.910 1140.670 ;
        RECT 1854.130 961.090 1855.310 962.270 ;
        RECT 1855.730 961.090 1856.910 962.270 ;
        RECT 1854.130 959.490 1855.310 960.670 ;
        RECT 1855.730 959.490 1856.910 960.670 ;
        RECT 1854.130 781.090 1855.310 782.270 ;
        RECT 1855.730 781.090 1856.910 782.270 ;
        RECT 1854.130 779.490 1855.310 780.670 ;
        RECT 1855.730 779.490 1856.910 780.670 ;
        RECT 1854.130 601.090 1855.310 602.270 ;
        RECT 1855.730 601.090 1856.910 602.270 ;
        RECT 1854.130 599.490 1855.310 600.670 ;
        RECT 1855.730 599.490 1856.910 600.670 ;
        RECT 1854.130 421.090 1855.310 422.270 ;
        RECT 1855.730 421.090 1856.910 422.270 ;
        RECT 1854.130 419.490 1855.310 420.670 ;
        RECT 1855.730 419.490 1856.910 420.670 ;
        RECT 1854.130 241.090 1855.310 242.270 ;
        RECT 1855.730 241.090 1856.910 242.270 ;
        RECT 1854.130 239.490 1855.310 240.670 ;
        RECT 1855.730 239.490 1856.910 240.670 ;
        RECT 1854.130 61.090 1855.310 62.270 ;
        RECT 1855.730 61.090 1856.910 62.270 ;
        RECT 1854.130 59.490 1855.310 60.670 ;
        RECT 1855.730 59.490 1856.910 60.670 ;
        RECT 1854.130 -12.510 1855.310 -11.330 ;
        RECT 1855.730 -12.510 1856.910 -11.330 ;
        RECT 1854.130 -14.110 1855.310 -12.930 ;
        RECT 1855.730 -14.110 1856.910 -12.930 ;
        RECT 2034.130 3532.610 2035.310 3533.790 ;
        RECT 2035.730 3532.610 2036.910 3533.790 ;
        RECT 2034.130 3531.010 2035.310 3532.190 ;
        RECT 2035.730 3531.010 2036.910 3532.190 ;
        RECT 2034.130 3481.090 2035.310 3482.270 ;
        RECT 2035.730 3481.090 2036.910 3482.270 ;
        RECT 2034.130 3479.490 2035.310 3480.670 ;
        RECT 2035.730 3479.490 2036.910 3480.670 ;
        RECT 2034.130 3301.090 2035.310 3302.270 ;
        RECT 2035.730 3301.090 2036.910 3302.270 ;
        RECT 2034.130 3299.490 2035.310 3300.670 ;
        RECT 2035.730 3299.490 2036.910 3300.670 ;
        RECT 2034.130 3121.090 2035.310 3122.270 ;
        RECT 2035.730 3121.090 2036.910 3122.270 ;
        RECT 2034.130 3119.490 2035.310 3120.670 ;
        RECT 2035.730 3119.490 2036.910 3120.670 ;
        RECT 2034.130 2941.090 2035.310 2942.270 ;
        RECT 2035.730 2941.090 2036.910 2942.270 ;
        RECT 2034.130 2939.490 2035.310 2940.670 ;
        RECT 2035.730 2939.490 2036.910 2940.670 ;
        RECT 2034.130 2761.090 2035.310 2762.270 ;
        RECT 2035.730 2761.090 2036.910 2762.270 ;
        RECT 2034.130 2759.490 2035.310 2760.670 ;
        RECT 2035.730 2759.490 2036.910 2760.670 ;
        RECT 2034.130 2581.090 2035.310 2582.270 ;
        RECT 2035.730 2581.090 2036.910 2582.270 ;
        RECT 2034.130 2579.490 2035.310 2580.670 ;
        RECT 2035.730 2579.490 2036.910 2580.670 ;
        RECT 2034.130 2401.090 2035.310 2402.270 ;
        RECT 2035.730 2401.090 2036.910 2402.270 ;
        RECT 2034.130 2399.490 2035.310 2400.670 ;
        RECT 2035.730 2399.490 2036.910 2400.670 ;
        RECT 2034.130 2221.090 2035.310 2222.270 ;
        RECT 2035.730 2221.090 2036.910 2222.270 ;
        RECT 2034.130 2219.490 2035.310 2220.670 ;
        RECT 2035.730 2219.490 2036.910 2220.670 ;
        RECT 2034.130 2041.090 2035.310 2042.270 ;
        RECT 2035.730 2041.090 2036.910 2042.270 ;
        RECT 2034.130 2039.490 2035.310 2040.670 ;
        RECT 2035.730 2039.490 2036.910 2040.670 ;
        RECT 2034.130 1861.090 2035.310 1862.270 ;
        RECT 2035.730 1861.090 2036.910 1862.270 ;
        RECT 2034.130 1859.490 2035.310 1860.670 ;
        RECT 2035.730 1859.490 2036.910 1860.670 ;
        RECT 2034.130 1681.090 2035.310 1682.270 ;
        RECT 2035.730 1681.090 2036.910 1682.270 ;
        RECT 2034.130 1679.490 2035.310 1680.670 ;
        RECT 2035.730 1679.490 2036.910 1680.670 ;
        RECT 2034.130 1501.090 2035.310 1502.270 ;
        RECT 2035.730 1501.090 2036.910 1502.270 ;
        RECT 2034.130 1499.490 2035.310 1500.670 ;
        RECT 2035.730 1499.490 2036.910 1500.670 ;
        RECT 2034.130 1321.090 2035.310 1322.270 ;
        RECT 2035.730 1321.090 2036.910 1322.270 ;
        RECT 2034.130 1319.490 2035.310 1320.670 ;
        RECT 2035.730 1319.490 2036.910 1320.670 ;
        RECT 2034.130 1141.090 2035.310 1142.270 ;
        RECT 2035.730 1141.090 2036.910 1142.270 ;
        RECT 2034.130 1139.490 2035.310 1140.670 ;
        RECT 2035.730 1139.490 2036.910 1140.670 ;
        RECT 2034.130 961.090 2035.310 962.270 ;
        RECT 2035.730 961.090 2036.910 962.270 ;
        RECT 2034.130 959.490 2035.310 960.670 ;
        RECT 2035.730 959.490 2036.910 960.670 ;
        RECT 2034.130 781.090 2035.310 782.270 ;
        RECT 2035.730 781.090 2036.910 782.270 ;
        RECT 2034.130 779.490 2035.310 780.670 ;
        RECT 2035.730 779.490 2036.910 780.670 ;
        RECT 2034.130 601.090 2035.310 602.270 ;
        RECT 2035.730 601.090 2036.910 602.270 ;
        RECT 2034.130 599.490 2035.310 600.670 ;
        RECT 2035.730 599.490 2036.910 600.670 ;
        RECT 2034.130 421.090 2035.310 422.270 ;
        RECT 2035.730 421.090 2036.910 422.270 ;
        RECT 2034.130 419.490 2035.310 420.670 ;
        RECT 2035.730 419.490 2036.910 420.670 ;
        RECT 2034.130 241.090 2035.310 242.270 ;
        RECT 2035.730 241.090 2036.910 242.270 ;
        RECT 2034.130 239.490 2035.310 240.670 ;
        RECT 2035.730 239.490 2036.910 240.670 ;
        RECT 2034.130 61.090 2035.310 62.270 ;
        RECT 2035.730 61.090 2036.910 62.270 ;
        RECT 2034.130 59.490 2035.310 60.670 ;
        RECT 2035.730 59.490 2036.910 60.670 ;
        RECT 2034.130 -12.510 2035.310 -11.330 ;
        RECT 2035.730 -12.510 2036.910 -11.330 ;
        RECT 2034.130 -14.110 2035.310 -12.930 ;
        RECT 2035.730 -14.110 2036.910 -12.930 ;
        RECT 2214.130 3532.610 2215.310 3533.790 ;
        RECT 2215.730 3532.610 2216.910 3533.790 ;
        RECT 2214.130 3531.010 2215.310 3532.190 ;
        RECT 2215.730 3531.010 2216.910 3532.190 ;
        RECT 2214.130 3481.090 2215.310 3482.270 ;
        RECT 2215.730 3481.090 2216.910 3482.270 ;
        RECT 2214.130 3479.490 2215.310 3480.670 ;
        RECT 2215.730 3479.490 2216.910 3480.670 ;
        RECT 2214.130 3301.090 2215.310 3302.270 ;
        RECT 2215.730 3301.090 2216.910 3302.270 ;
        RECT 2214.130 3299.490 2215.310 3300.670 ;
        RECT 2215.730 3299.490 2216.910 3300.670 ;
        RECT 2214.130 3121.090 2215.310 3122.270 ;
        RECT 2215.730 3121.090 2216.910 3122.270 ;
        RECT 2214.130 3119.490 2215.310 3120.670 ;
        RECT 2215.730 3119.490 2216.910 3120.670 ;
        RECT 2214.130 2941.090 2215.310 2942.270 ;
        RECT 2215.730 2941.090 2216.910 2942.270 ;
        RECT 2214.130 2939.490 2215.310 2940.670 ;
        RECT 2215.730 2939.490 2216.910 2940.670 ;
        RECT 2214.130 2761.090 2215.310 2762.270 ;
        RECT 2215.730 2761.090 2216.910 2762.270 ;
        RECT 2214.130 2759.490 2215.310 2760.670 ;
        RECT 2215.730 2759.490 2216.910 2760.670 ;
        RECT 2214.130 2581.090 2215.310 2582.270 ;
        RECT 2215.730 2581.090 2216.910 2582.270 ;
        RECT 2214.130 2579.490 2215.310 2580.670 ;
        RECT 2215.730 2579.490 2216.910 2580.670 ;
        RECT 2214.130 2401.090 2215.310 2402.270 ;
        RECT 2215.730 2401.090 2216.910 2402.270 ;
        RECT 2214.130 2399.490 2215.310 2400.670 ;
        RECT 2215.730 2399.490 2216.910 2400.670 ;
        RECT 2214.130 2221.090 2215.310 2222.270 ;
        RECT 2215.730 2221.090 2216.910 2222.270 ;
        RECT 2214.130 2219.490 2215.310 2220.670 ;
        RECT 2215.730 2219.490 2216.910 2220.670 ;
        RECT 2214.130 2041.090 2215.310 2042.270 ;
        RECT 2215.730 2041.090 2216.910 2042.270 ;
        RECT 2214.130 2039.490 2215.310 2040.670 ;
        RECT 2215.730 2039.490 2216.910 2040.670 ;
        RECT 2214.130 1861.090 2215.310 1862.270 ;
        RECT 2215.730 1861.090 2216.910 1862.270 ;
        RECT 2214.130 1859.490 2215.310 1860.670 ;
        RECT 2215.730 1859.490 2216.910 1860.670 ;
        RECT 2214.130 1681.090 2215.310 1682.270 ;
        RECT 2215.730 1681.090 2216.910 1682.270 ;
        RECT 2214.130 1679.490 2215.310 1680.670 ;
        RECT 2215.730 1679.490 2216.910 1680.670 ;
        RECT 2214.130 1501.090 2215.310 1502.270 ;
        RECT 2215.730 1501.090 2216.910 1502.270 ;
        RECT 2214.130 1499.490 2215.310 1500.670 ;
        RECT 2215.730 1499.490 2216.910 1500.670 ;
        RECT 2214.130 1321.090 2215.310 1322.270 ;
        RECT 2215.730 1321.090 2216.910 1322.270 ;
        RECT 2214.130 1319.490 2215.310 1320.670 ;
        RECT 2215.730 1319.490 2216.910 1320.670 ;
        RECT 2214.130 1141.090 2215.310 1142.270 ;
        RECT 2215.730 1141.090 2216.910 1142.270 ;
        RECT 2214.130 1139.490 2215.310 1140.670 ;
        RECT 2215.730 1139.490 2216.910 1140.670 ;
        RECT 2214.130 961.090 2215.310 962.270 ;
        RECT 2215.730 961.090 2216.910 962.270 ;
        RECT 2214.130 959.490 2215.310 960.670 ;
        RECT 2215.730 959.490 2216.910 960.670 ;
        RECT 2214.130 781.090 2215.310 782.270 ;
        RECT 2215.730 781.090 2216.910 782.270 ;
        RECT 2214.130 779.490 2215.310 780.670 ;
        RECT 2215.730 779.490 2216.910 780.670 ;
        RECT 2214.130 601.090 2215.310 602.270 ;
        RECT 2215.730 601.090 2216.910 602.270 ;
        RECT 2214.130 599.490 2215.310 600.670 ;
        RECT 2215.730 599.490 2216.910 600.670 ;
        RECT 2214.130 421.090 2215.310 422.270 ;
        RECT 2215.730 421.090 2216.910 422.270 ;
        RECT 2214.130 419.490 2215.310 420.670 ;
        RECT 2215.730 419.490 2216.910 420.670 ;
        RECT 2214.130 241.090 2215.310 242.270 ;
        RECT 2215.730 241.090 2216.910 242.270 ;
        RECT 2214.130 239.490 2215.310 240.670 ;
        RECT 2215.730 239.490 2216.910 240.670 ;
        RECT 2214.130 61.090 2215.310 62.270 ;
        RECT 2215.730 61.090 2216.910 62.270 ;
        RECT 2214.130 59.490 2215.310 60.670 ;
        RECT 2215.730 59.490 2216.910 60.670 ;
        RECT 2214.130 -12.510 2215.310 -11.330 ;
        RECT 2215.730 -12.510 2216.910 -11.330 ;
        RECT 2214.130 -14.110 2215.310 -12.930 ;
        RECT 2215.730 -14.110 2216.910 -12.930 ;
        RECT 2394.130 3532.610 2395.310 3533.790 ;
        RECT 2395.730 3532.610 2396.910 3533.790 ;
        RECT 2394.130 3531.010 2395.310 3532.190 ;
        RECT 2395.730 3531.010 2396.910 3532.190 ;
        RECT 2394.130 3481.090 2395.310 3482.270 ;
        RECT 2395.730 3481.090 2396.910 3482.270 ;
        RECT 2394.130 3479.490 2395.310 3480.670 ;
        RECT 2395.730 3479.490 2396.910 3480.670 ;
        RECT 2394.130 3301.090 2395.310 3302.270 ;
        RECT 2395.730 3301.090 2396.910 3302.270 ;
        RECT 2394.130 3299.490 2395.310 3300.670 ;
        RECT 2395.730 3299.490 2396.910 3300.670 ;
        RECT 2394.130 3121.090 2395.310 3122.270 ;
        RECT 2395.730 3121.090 2396.910 3122.270 ;
        RECT 2394.130 3119.490 2395.310 3120.670 ;
        RECT 2395.730 3119.490 2396.910 3120.670 ;
        RECT 2394.130 2941.090 2395.310 2942.270 ;
        RECT 2395.730 2941.090 2396.910 2942.270 ;
        RECT 2394.130 2939.490 2395.310 2940.670 ;
        RECT 2395.730 2939.490 2396.910 2940.670 ;
        RECT 2394.130 2761.090 2395.310 2762.270 ;
        RECT 2395.730 2761.090 2396.910 2762.270 ;
        RECT 2394.130 2759.490 2395.310 2760.670 ;
        RECT 2395.730 2759.490 2396.910 2760.670 ;
        RECT 2394.130 2581.090 2395.310 2582.270 ;
        RECT 2395.730 2581.090 2396.910 2582.270 ;
        RECT 2394.130 2579.490 2395.310 2580.670 ;
        RECT 2395.730 2579.490 2396.910 2580.670 ;
        RECT 2394.130 2401.090 2395.310 2402.270 ;
        RECT 2395.730 2401.090 2396.910 2402.270 ;
        RECT 2394.130 2399.490 2395.310 2400.670 ;
        RECT 2395.730 2399.490 2396.910 2400.670 ;
        RECT 2394.130 2221.090 2395.310 2222.270 ;
        RECT 2395.730 2221.090 2396.910 2222.270 ;
        RECT 2394.130 2219.490 2395.310 2220.670 ;
        RECT 2395.730 2219.490 2396.910 2220.670 ;
        RECT 2394.130 2041.090 2395.310 2042.270 ;
        RECT 2395.730 2041.090 2396.910 2042.270 ;
        RECT 2394.130 2039.490 2395.310 2040.670 ;
        RECT 2395.730 2039.490 2396.910 2040.670 ;
        RECT 2394.130 1861.090 2395.310 1862.270 ;
        RECT 2395.730 1861.090 2396.910 1862.270 ;
        RECT 2394.130 1859.490 2395.310 1860.670 ;
        RECT 2395.730 1859.490 2396.910 1860.670 ;
        RECT 2394.130 1681.090 2395.310 1682.270 ;
        RECT 2395.730 1681.090 2396.910 1682.270 ;
        RECT 2394.130 1679.490 2395.310 1680.670 ;
        RECT 2395.730 1679.490 2396.910 1680.670 ;
        RECT 2394.130 1501.090 2395.310 1502.270 ;
        RECT 2395.730 1501.090 2396.910 1502.270 ;
        RECT 2394.130 1499.490 2395.310 1500.670 ;
        RECT 2395.730 1499.490 2396.910 1500.670 ;
        RECT 2394.130 1321.090 2395.310 1322.270 ;
        RECT 2395.730 1321.090 2396.910 1322.270 ;
        RECT 2394.130 1319.490 2395.310 1320.670 ;
        RECT 2395.730 1319.490 2396.910 1320.670 ;
        RECT 2394.130 1141.090 2395.310 1142.270 ;
        RECT 2395.730 1141.090 2396.910 1142.270 ;
        RECT 2394.130 1139.490 2395.310 1140.670 ;
        RECT 2395.730 1139.490 2396.910 1140.670 ;
        RECT 2394.130 961.090 2395.310 962.270 ;
        RECT 2395.730 961.090 2396.910 962.270 ;
        RECT 2394.130 959.490 2395.310 960.670 ;
        RECT 2395.730 959.490 2396.910 960.670 ;
        RECT 2394.130 781.090 2395.310 782.270 ;
        RECT 2395.730 781.090 2396.910 782.270 ;
        RECT 2394.130 779.490 2395.310 780.670 ;
        RECT 2395.730 779.490 2396.910 780.670 ;
        RECT 2394.130 601.090 2395.310 602.270 ;
        RECT 2395.730 601.090 2396.910 602.270 ;
        RECT 2394.130 599.490 2395.310 600.670 ;
        RECT 2395.730 599.490 2396.910 600.670 ;
        RECT 2394.130 421.090 2395.310 422.270 ;
        RECT 2395.730 421.090 2396.910 422.270 ;
        RECT 2394.130 419.490 2395.310 420.670 ;
        RECT 2395.730 419.490 2396.910 420.670 ;
        RECT 2394.130 241.090 2395.310 242.270 ;
        RECT 2395.730 241.090 2396.910 242.270 ;
        RECT 2394.130 239.490 2395.310 240.670 ;
        RECT 2395.730 239.490 2396.910 240.670 ;
        RECT 2394.130 61.090 2395.310 62.270 ;
        RECT 2395.730 61.090 2396.910 62.270 ;
        RECT 2394.130 59.490 2395.310 60.670 ;
        RECT 2395.730 59.490 2396.910 60.670 ;
        RECT 2394.130 -12.510 2395.310 -11.330 ;
        RECT 2395.730 -12.510 2396.910 -11.330 ;
        RECT 2394.130 -14.110 2395.310 -12.930 ;
        RECT 2395.730 -14.110 2396.910 -12.930 ;
        RECT 2574.130 3532.610 2575.310 3533.790 ;
        RECT 2575.730 3532.610 2576.910 3533.790 ;
        RECT 2574.130 3531.010 2575.310 3532.190 ;
        RECT 2575.730 3531.010 2576.910 3532.190 ;
        RECT 2574.130 3481.090 2575.310 3482.270 ;
        RECT 2575.730 3481.090 2576.910 3482.270 ;
        RECT 2574.130 3479.490 2575.310 3480.670 ;
        RECT 2575.730 3479.490 2576.910 3480.670 ;
        RECT 2574.130 3301.090 2575.310 3302.270 ;
        RECT 2575.730 3301.090 2576.910 3302.270 ;
        RECT 2574.130 3299.490 2575.310 3300.670 ;
        RECT 2575.730 3299.490 2576.910 3300.670 ;
        RECT 2574.130 3121.090 2575.310 3122.270 ;
        RECT 2575.730 3121.090 2576.910 3122.270 ;
        RECT 2574.130 3119.490 2575.310 3120.670 ;
        RECT 2575.730 3119.490 2576.910 3120.670 ;
        RECT 2574.130 2941.090 2575.310 2942.270 ;
        RECT 2575.730 2941.090 2576.910 2942.270 ;
        RECT 2574.130 2939.490 2575.310 2940.670 ;
        RECT 2575.730 2939.490 2576.910 2940.670 ;
        RECT 2574.130 2761.090 2575.310 2762.270 ;
        RECT 2575.730 2761.090 2576.910 2762.270 ;
        RECT 2574.130 2759.490 2575.310 2760.670 ;
        RECT 2575.730 2759.490 2576.910 2760.670 ;
        RECT 2574.130 2581.090 2575.310 2582.270 ;
        RECT 2575.730 2581.090 2576.910 2582.270 ;
        RECT 2574.130 2579.490 2575.310 2580.670 ;
        RECT 2575.730 2579.490 2576.910 2580.670 ;
        RECT 2574.130 2401.090 2575.310 2402.270 ;
        RECT 2575.730 2401.090 2576.910 2402.270 ;
        RECT 2574.130 2399.490 2575.310 2400.670 ;
        RECT 2575.730 2399.490 2576.910 2400.670 ;
        RECT 2574.130 2221.090 2575.310 2222.270 ;
        RECT 2575.730 2221.090 2576.910 2222.270 ;
        RECT 2574.130 2219.490 2575.310 2220.670 ;
        RECT 2575.730 2219.490 2576.910 2220.670 ;
        RECT 2574.130 2041.090 2575.310 2042.270 ;
        RECT 2575.730 2041.090 2576.910 2042.270 ;
        RECT 2574.130 2039.490 2575.310 2040.670 ;
        RECT 2575.730 2039.490 2576.910 2040.670 ;
        RECT 2574.130 1861.090 2575.310 1862.270 ;
        RECT 2575.730 1861.090 2576.910 1862.270 ;
        RECT 2574.130 1859.490 2575.310 1860.670 ;
        RECT 2575.730 1859.490 2576.910 1860.670 ;
        RECT 2574.130 1681.090 2575.310 1682.270 ;
        RECT 2575.730 1681.090 2576.910 1682.270 ;
        RECT 2574.130 1679.490 2575.310 1680.670 ;
        RECT 2575.730 1679.490 2576.910 1680.670 ;
        RECT 2574.130 1501.090 2575.310 1502.270 ;
        RECT 2575.730 1501.090 2576.910 1502.270 ;
        RECT 2574.130 1499.490 2575.310 1500.670 ;
        RECT 2575.730 1499.490 2576.910 1500.670 ;
        RECT 2574.130 1321.090 2575.310 1322.270 ;
        RECT 2575.730 1321.090 2576.910 1322.270 ;
        RECT 2574.130 1319.490 2575.310 1320.670 ;
        RECT 2575.730 1319.490 2576.910 1320.670 ;
        RECT 2574.130 1141.090 2575.310 1142.270 ;
        RECT 2575.730 1141.090 2576.910 1142.270 ;
        RECT 2574.130 1139.490 2575.310 1140.670 ;
        RECT 2575.730 1139.490 2576.910 1140.670 ;
        RECT 2574.130 961.090 2575.310 962.270 ;
        RECT 2575.730 961.090 2576.910 962.270 ;
        RECT 2574.130 959.490 2575.310 960.670 ;
        RECT 2575.730 959.490 2576.910 960.670 ;
        RECT 2574.130 781.090 2575.310 782.270 ;
        RECT 2575.730 781.090 2576.910 782.270 ;
        RECT 2574.130 779.490 2575.310 780.670 ;
        RECT 2575.730 779.490 2576.910 780.670 ;
        RECT 2574.130 601.090 2575.310 602.270 ;
        RECT 2575.730 601.090 2576.910 602.270 ;
        RECT 2574.130 599.490 2575.310 600.670 ;
        RECT 2575.730 599.490 2576.910 600.670 ;
        RECT 2574.130 421.090 2575.310 422.270 ;
        RECT 2575.730 421.090 2576.910 422.270 ;
        RECT 2574.130 419.490 2575.310 420.670 ;
        RECT 2575.730 419.490 2576.910 420.670 ;
        RECT 2574.130 241.090 2575.310 242.270 ;
        RECT 2575.730 241.090 2576.910 242.270 ;
        RECT 2574.130 239.490 2575.310 240.670 ;
        RECT 2575.730 239.490 2576.910 240.670 ;
        RECT 2574.130 61.090 2575.310 62.270 ;
        RECT 2575.730 61.090 2576.910 62.270 ;
        RECT 2574.130 59.490 2575.310 60.670 ;
        RECT 2575.730 59.490 2576.910 60.670 ;
        RECT 2574.130 -12.510 2575.310 -11.330 ;
        RECT 2575.730 -12.510 2576.910 -11.330 ;
        RECT 2574.130 -14.110 2575.310 -12.930 ;
        RECT 2575.730 -14.110 2576.910 -12.930 ;
        RECT 2754.130 3532.610 2755.310 3533.790 ;
        RECT 2755.730 3532.610 2756.910 3533.790 ;
        RECT 2754.130 3531.010 2755.310 3532.190 ;
        RECT 2755.730 3531.010 2756.910 3532.190 ;
        RECT 2754.130 3481.090 2755.310 3482.270 ;
        RECT 2755.730 3481.090 2756.910 3482.270 ;
        RECT 2754.130 3479.490 2755.310 3480.670 ;
        RECT 2755.730 3479.490 2756.910 3480.670 ;
        RECT 2754.130 3301.090 2755.310 3302.270 ;
        RECT 2755.730 3301.090 2756.910 3302.270 ;
        RECT 2754.130 3299.490 2755.310 3300.670 ;
        RECT 2755.730 3299.490 2756.910 3300.670 ;
        RECT 2754.130 3121.090 2755.310 3122.270 ;
        RECT 2755.730 3121.090 2756.910 3122.270 ;
        RECT 2754.130 3119.490 2755.310 3120.670 ;
        RECT 2755.730 3119.490 2756.910 3120.670 ;
        RECT 2754.130 2941.090 2755.310 2942.270 ;
        RECT 2755.730 2941.090 2756.910 2942.270 ;
        RECT 2754.130 2939.490 2755.310 2940.670 ;
        RECT 2755.730 2939.490 2756.910 2940.670 ;
        RECT 2754.130 2761.090 2755.310 2762.270 ;
        RECT 2755.730 2761.090 2756.910 2762.270 ;
        RECT 2754.130 2759.490 2755.310 2760.670 ;
        RECT 2755.730 2759.490 2756.910 2760.670 ;
        RECT 2754.130 2581.090 2755.310 2582.270 ;
        RECT 2755.730 2581.090 2756.910 2582.270 ;
        RECT 2754.130 2579.490 2755.310 2580.670 ;
        RECT 2755.730 2579.490 2756.910 2580.670 ;
        RECT 2754.130 2401.090 2755.310 2402.270 ;
        RECT 2755.730 2401.090 2756.910 2402.270 ;
        RECT 2754.130 2399.490 2755.310 2400.670 ;
        RECT 2755.730 2399.490 2756.910 2400.670 ;
        RECT 2754.130 2221.090 2755.310 2222.270 ;
        RECT 2755.730 2221.090 2756.910 2222.270 ;
        RECT 2754.130 2219.490 2755.310 2220.670 ;
        RECT 2755.730 2219.490 2756.910 2220.670 ;
        RECT 2754.130 2041.090 2755.310 2042.270 ;
        RECT 2755.730 2041.090 2756.910 2042.270 ;
        RECT 2754.130 2039.490 2755.310 2040.670 ;
        RECT 2755.730 2039.490 2756.910 2040.670 ;
        RECT 2754.130 1861.090 2755.310 1862.270 ;
        RECT 2755.730 1861.090 2756.910 1862.270 ;
        RECT 2754.130 1859.490 2755.310 1860.670 ;
        RECT 2755.730 1859.490 2756.910 1860.670 ;
        RECT 2754.130 1681.090 2755.310 1682.270 ;
        RECT 2755.730 1681.090 2756.910 1682.270 ;
        RECT 2754.130 1679.490 2755.310 1680.670 ;
        RECT 2755.730 1679.490 2756.910 1680.670 ;
        RECT 2754.130 1501.090 2755.310 1502.270 ;
        RECT 2755.730 1501.090 2756.910 1502.270 ;
        RECT 2754.130 1499.490 2755.310 1500.670 ;
        RECT 2755.730 1499.490 2756.910 1500.670 ;
        RECT 2754.130 1321.090 2755.310 1322.270 ;
        RECT 2755.730 1321.090 2756.910 1322.270 ;
        RECT 2754.130 1319.490 2755.310 1320.670 ;
        RECT 2755.730 1319.490 2756.910 1320.670 ;
        RECT 2754.130 1141.090 2755.310 1142.270 ;
        RECT 2755.730 1141.090 2756.910 1142.270 ;
        RECT 2754.130 1139.490 2755.310 1140.670 ;
        RECT 2755.730 1139.490 2756.910 1140.670 ;
        RECT 2754.130 961.090 2755.310 962.270 ;
        RECT 2755.730 961.090 2756.910 962.270 ;
        RECT 2754.130 959.490 2755.310 960.670 ;
        RECT 2755.730 959.490 2756.910 960.670 ;
        RECT 2754.130 781.090 2755.310 782.270 ;
        RECT 2755.730 781.090 2756.910 782.270 ;
        RECT 2754.130 779.490 2755.310 780.670 ;
        RECT 2755.730 779.490 2756.910 780.670 ;
        RECT 2754.130 601.090 2755.310 602.270 ;
        RECT 2755.730 601.090 2756.910 602.270 ;
        RECT 2754.130 599.490 2755.310 600.670 ;
        RECT 2755.730 599.490 2756.910 600.670 ;
        RECT 2754.130 421.090 2755.310 422.270 ;
        RECT 2755.730 421.090 2756.910 422.270 ;
        RECT 2754.130 419.490 2755.310 420.670 ;
        RECT 2755.730 419.490 2756.910 420.670 ;
        RECT 2754.130 241.090 2755.310 242.270 ;
        RECT 2755.730 241.090 2756.910 242.270 ;
        RECT 2754.130 239.490 2755.310 240.670 ;
        RECT 2755.730 239.490 2756.910 240.670 ;
        RECT 2754.130 61.090 2755.310 62.270 ;
        RECT 2755.730 61.090 2756.910 62.270 ;
        RECT 2754.130 59.490 2755.310 60.670 ;
        RECT 2755.730 59.490 2756.910 60.670 ;
        RECT 2754.130 -12.510 2755.310 -11.330 ;
        RECT 2755.730 -12.510 2756.910 -11.330 ;
        RECT 2754.130 -14.110 2755.310 -12.930 ;
        RECT 2755.730 -14.110 2756.910 -12.930 ;
        RECT 2936.310 3532.610 2937.490 3533.790 ;
        RECT 2937.910 3532.610 2939.090 3533.790 ;
        RECT 2936.310 3531.010 2937.490 3532.190 ;
        RECT 2937.910 3531.010 2939.090 3532.190 ;
        RECT 2936.310 3481.090 2937.490 3482.270 ;
        RECT 2937.910 3481.090 2939.090 3482.270 ;
        RECT 2936.310 3479.490 2937.490 3480.670 ;
        RECT 2937.910 3479.490 2939.090 3480.670 ;
        RECT 2936.310 3301.090 2937.490 3302.270 ;
        RECT 2937.910 3301.090 2939.090 3302.270 ;
        RECT 2936.310 3299.490 2937.490 3300.670 ;
        RECT 2937.910 3299.490 2939.090 3300.670 ;
        RECT 2936.310 3121.090 2937.490 3122.270 ;
        RECT 2937.910 3121.090 2939.090 3122.270 ;
        RECT 2936.310 3119.490 2937.490 3120.670 ;
        RECT 2937.910 3119.490 2939.090 3120.670 ;
        RECT 2936.310 2941.090 2937.490 2942.270 ;
        RECT 2937.910 2941.090 2939.090 2942.270 ;
        RECT 2936.310 2939.490 2937.490 2940.670 ;
        RECT 2937.910 2939.490 2939.090 2940.670 ;
        RECT 2936.310 2761.090 2937.490 2762.270 ;
        RECT 2937.910 2761.090 2939.090 2762.270 ;
        RECT 2936.310 2759.490 2937.490 2760.670 ;
        RECT 2937.910 2759.490 2939.090 2760.670 ;
        RECT 2936.310 2581.090 2937.490 2582.270 ;
        RECT 2937.910 2581.090 2939.090 2582.270 ;
        RECT 2936.310 2579.490 2937.490 2580.670 ;
        RECT 2937.910 2579.490 2939.090 2580.670 ;
        RECT 2936.310 2401.090 2937.490 2402.270 ;
        RECT 2937.910 2401.090 2939.090 2402.270 ;
        RECT 2936.310 2399.490 2937.490 2400.670 ;
        RECT 2937.910 2399.490 2939.090 2400.670 ;
        RECT 2936.310 2221.090 2937.490 2222.270 ;
        RECT 2937.910 2221.090 2939.090 2222.270 ;
        RECT 2936.310 2219.490 2937.490 2220.670 ;
        RECT 2937.910 2219.490 2939.090 2220.670 ;
        RECT 2936.310 2041.090 2937.490 2042.270 ;
        RECT 2937.910 2041.090 2939.090 2042.270 ;
        RECT 2936.310 2039.490 2937.490 2040.670 ;
        RECT 2937.910 2039.490 2939.090 2040.670 ;
        RECT 2936.310 1861.090 2937.490 1862.270 ;
        RECT 2937.910 1861.090 2939.090 1862.270 ;
        RECT 2936.310 1859.490 2937.490 1860.670 ;
        RECT 2937.910 1859.490 2939.090 1860.670 ;
        RECT 2936.310 1681.090 2937.490 1682.270 ;
        RECT 2937.910 1681.090 2939.090 1682.270 ;
        RECT 2936.310 1679.490 2937.490 1680.670 ;
        RECT 2937.910 1679.490 2939.090 1680.670 ;
        RECT 2936.310 1501.090 2937.490 1502.270 ;
        RECT 2937.910 1501.090 2939.090 1502.270 ;
        RECT 2936.310 1499.490 2937.490 1500.670 ;
        RECT 2937.910 1499.490 2939.090 1500.670 ;
        RECT 2936.310 1321.090 2937.490 1322.270 ;
        RECT 2937.910 1321.090 2939.090 1322.270 ;
        RECT 2936.310 1319.490 2937.490 1320.670 ;
        RECT 2937.910 1319.490 2939.090 1320.670 ;
        RECT 2936.310 1141.090 2937.490 1142.270 ;
        RECT 2937.910 1141.090 2939.090 1142.270 ;
        RECT 2936.310 1139.490 2937.490 1140.670 ;
        RECT 2937.910 1139.490 2939.090 1140.670 ;
        RECT 2936.310 961.090 2937.490 962.270 ;
        RECT 2937.910 961.090 2939.090 962.270 ;
        RECT 2936.310 959.490 2937.490 960.670 ;
        RECT 2937.910 959.490 2939.090 960.670 ;
        RECT 2936.310 781.090 2937.490 782.270 ;
        RECT 2937.910 781.090 2939.090 782.270 ;
        RECT 2936.310 779.490 2937.490 780.670 ;
        RECT 2937.910 779.490 2939.090 780.670 ;
        RECT 2936.310 601.090 2937.490 602.270 ;
        RECT 2937.910 601.090 2939.090 602.270 ;
        RECT 2936.310 599.490 2937.490 600.670 ;
        RECT 2937.910 599.490 2939.090 600.670 ;
        RECT 2936.310 421.090 2937.490 422.270 ;
        RECT 2937.910 421.090 2939.090 422.270 ;
        RECT 2936.310 419.490 2937.490 420.670 ;
        RECT 2937.910 419.490 2939.090 420.670 ;
        RECT 2936.310 241.090 2937.490 242.270 ;
        RECT 2937.910 241.090 2939.090 242.270 ;
        RECT 2936.310 239.490 2937.490 240.670 ;
        RECT 2937.910 239.490 2939.090 240.670 ;
        RECT 2936.310 61.090 2937.490 62.270 ;
        RECT 2937.910 61.090 2939.090 62.270 ;
        RECT 2936.310 59.490 2937.490 60.670 ;
        RECT 2937.910 59.490 2939.090 60.670 ;
        RECT 2936.310 -12.510 2937.490 -11.330 ;
        RECT 2937.910 -12.510 2939.090 -11.330 ;
        RECT 2936.310 -14.110 2937.490 -12.930 ;
        RECT 2937.910 -14.110 2939.090 -12.930 ;
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
        RECT -43.630 3479.330 2963.250 3482.430 ;
        RECT -43.630 3299.330 2963.250 3302.430 ;
        RECT -43.630 3119.330 2963.250 3122.430 ;
        RECT -43.630 2939.330 2963.250 2942.430 ;
        RECT -43.630 2759.330 2963.250 2762.430 ;
        RECT -43.630 2579.330 2963.250 2582.430 ;
        RECT -43.630 2399.330 2963.250 2402.430 ;
        RECT -43.630 2219.330 2963.250 2222.430 ;
        RECT -43.630 2039.330 2963.250 2042.430 ;
        RECT -43.630 1859.330 2963.250 1862.430 ;
        RECT -43.630 1679.330 2963.250 1682.430 ;
        RECT -43.630 1499.330 2963.250 1502.430 ;
        RECT -43.630 1319.330 2963.250 1322.430 ;
        RECT -43.630 1139.330 2963.250 1142.430 ;
        RECT -43.630 959.330 2963.250 962.430 ;
        RECT -43.630 779.330 2963.250 782.430 ;
        RECT -43.630 599.330 2963.250 602.430 ;
        RECT -43.630 419.330 2963.250 422.430 ;
        RECT -43.630 239.330 2963.250 242.430 ;
        RECT -43.630 59.330 2963.250 62.430 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
        RECT 98.970 -38.270 102.070 3557.950 ;
        RECT 278.970 -38.270 282.070 3557.950 ;
        RECT 458.970 810.000 462.070 3557.950 ;
        RECT 638.970 810.000 642.070 3557.950 ;
        RECT 458.970 -38.270 462.070 490.000 ;
        RECT 638.970 -38.270 642.070 490.000 ;
        RECT 818.970 -38.270 822.070 3557.950 ;
        RECT 998.970 -38.270 1002.070 3557.950 ;
        RECT 1178.970 -38.270 1182.070 3557.950 ;
        RECT 1358.970 -38.270 1362.070 3557.950 ;
        RECT 1538.970 -38.270 1542.070 3557.950 ;
        RECT 1718.970 -38.270 1722.070 3557.950 ;
        RECT 1898.970 -38.270 1902.070 3557.950 ;
        RECT 2078.970 -38.270 2082.070 3557.950 ;
        RECT 2258.970 -38.270 2262.070 3557.950 ;
        RECT 2438.970 -38.270 2442.070 3557.950 ;
        RECT 2618.970 -38.270 2622.070 3557.950 ;
        RECT 2798.970 -38.270 2802.070 3557.950 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
      LAYER via4 ;
        RECT -29.070 3542.210 -27.890 3543.390 ;
        RECT -27.470 3542.210 -26.290 3543.390 ;
        RECT -29.070 3540.610 -27.890 3541.790 ;
        RECT -27.470 3540.610 -26.290 3541.790 ;
        RECT -29.070 3346.090 -27.890 3347.270 ;
        RECT -27.470 3346.090 -26.290 3347.270 ;
        RECT -29.070 3344.490 -27.890 3345.670 ;
        RECT -27.470 3344.490 -26.290 3345.670 ;
        RECT -29.070 3166.090 -27.890 3167.270 ;
        RECT -27.470 3166.090 -26.290 3167.270 ;
        RECT -29.070 3164.490 -27.890 3165.670 ;
        RECT -27.470 3164.490 -26.290 3165.670 ;
        RECT -29.070 2986.090 -27.890 2987.270 ;
        RECT -27.470 2986.090 -26.290 2987.270 ;
        RECT -29.070 2984.490 -27.890 2985.670 ;
        RECT -27.470 2984.490 -26.290 2985.670 ;
        RECT -29.070 2806.090 -27.890 2807.270 ;
        RECT -27.470 2806.090 -26.290 2807.270 ;
        RECT -29.070 2804.490 -27.890 2805.670 ;
        RECT -27.470 2804.490 -26.290 2805.670 ;
        RECT -29.070 2626.090 -27.890 2627.270 ;
        RECT -27.470 2626.090 -26.290 2627.270 ;
        RECT -29.070 2624.490 -27.890 2625.670 ;
        RECT -27.470 2624.490 -26.290 2625.670 ;
        RECT -29.070 2446.090 -27.890 2447.270 ;
        RECT -27.470 2446.090 -26.290 2447.270 ;
        RECT -29.070 2444.490 -27.890 2445.670 ;
        RECT -27.470 2444.490 -26.290 2445.670 ;
        RECT -29.070 2266.090 -27.890 2267.270 ;
        RECT -27.470 2266.090 -26.290 2267.270 ;
        RECT -29.070 2264.490 -27.890 2265.670 ;
        RECT -27.470 2264.490 -26.290 2265.670 ;
        RECT -29.070 2086.090 -27.890 2087.270 ;
        RECT -27.470 2086.090 -26.290 2087.270 ;
        RECT -29.070 2084.490 -27.890 2085.670 ;
        RECT -27.470 2084.490 -26.290 2085.670 ;
        RECT -29.070 1906.090 -27.890 1907.270 ;
        RECT -27.470 1906.090 -26.290 1907.270 ;
        RECT -29.070 1904.490 -27.890 1905.670 ;
        RECT -27.470 1904.490 -26.290 1905.670 ;
        RECT -29.070 1726.090 -27.890 1727.270 ;
        RECT -27.470 1726.090 -26.290 1727.270 ;
        RECT -29.070 1724.490 -27.890 1725.670 ;
        RECT -27.470 1724.490 -26.290 1725.670 ;
        RECT -29.070 1546.090 -27.890 1547.270 ;
        RECT -27.470 1546.090 -26.290 1547.270 ;
        RECT -29.070 1544.490 -27.890 1545.670 ;
        RECT -27.470 1544.490 -26.290 1545.670 ;
        RECT -29.070 1366.090 -27.890 1367.270 ;
        RECT -27.470 1366.090 -26.290 1367.270 ;
        RECT -29.070 1364.490 -27.890 1365.670 ;
        RECT -27.470 1364.490 -26.290 1365.670 ;
        RECT -29.070 1186.090 -27.890 1187.270 ;
        RECT -27.470 1186.090 -26.290 1187.270 ;
        RECT -29.070 1184.490 -27.890 1185.670 ;
        RECT -27.470 1184.490 -26.290 1185.670 ;
        RECT -29.070 1006.090 -27.890 1007.270 ;
        RECT -27.470 1006.090 -26.290 1007.270 ;
        RECT -29.070 1004.490 -27.890 1005.670 ;
        RECT -27.470 1004.490 -26.290 1005.670 ;
        RECT -29.070 826.090 -27.890 827.270 ;
        RECT -27.470 826.090 -26.290 827.270 ;
        RECT -29.070 824.490 -27.890 825.670 ;
        RECT -27.470 824.490 -26.290 825.670 ;
        RECT -29.070 646.090 -27.890 647.270 ;
        RECT -27.470 646.090 -26.290 647.270 ;
        RECT -29.070 644.490 -27.890 645.670 ;
        RECT -27.470 644.490 -26.290 645.670 ;
        RECT -29.070 466.090 -27.890 467.270 ;
        RECT -27.470 466.090 -26.290 467.270 ;
        RECT -29.070 464.490 -27.890 465.670 ;
        RECT -27.470 464.490 -26.290 465.670 ;
        RECT -29.070 286.090 -27.890 287.270 ;
        RECT -27.470 286.090 -26.290 287.270 ;
        RECT -29.070 284.490 -27.890 285.670 ;
        RECT -27.470 284.490 -26.290 285.670 ;
        RECT -29.070 106.090 -27.890 107.270 ;
        RECT -27.470 106.090 -26.290 107.270 ;
        RECT -29.070 104.490 -27.890 105.670 ;
        RECT -27.470 104.490 -26.290 105.670 ;
        RECT -29.070 -22.110 -27.890 -20.930 ;
        RECT -27.470 -22.110 -26.290 -20.930 ;
        RECT -29.070 -23.710 -27.890 -22.530 ;
        RECT -27.470 -23.710 -26.290 -22.530 ;
        RECT 99.130 3542.210 100.310 3543.390 ;
        RECT 100.730 3542.210 101.910 3543.390 ;
        RECT 99.130 3540.610 100.310 3541.790 ;
        RECT 100.730 3540.610 101.910 3541.790 ;
        RECT 99.130 3346.090 100.310 3347.270 ;
        RECT 100.730 3346.090 101.910 3347.270 ;
        RECT 99.130 3344.490 100.310 3345.670 ;
        RECT 100.730 3344.490 101.910 3345.670 ;
        RECT 99.130 3166.090 100.310 3167.270 ;
        RECT 100.730 3166.090 101.910 3167.270 ;
        RECT 99.130 3164.490 100.310 3165.670 ;
        RECT 100.730 3164.490 101.910 3165.670 ;
        RECT 99.130 2986.090 100.310 2987.270 ;
        RECT 100.730 2986.090 101.910 2987.270 ;
        RECT 99.130 2984.490 100.310 2985.670 ;
        RECT 100.730 2984.490 101.910 2985.670 ;
        RECT 99.130 2806.090 100.310 2807.270 ;
        RECT 100.730 2806.090 101.910 2807.270 ;
        RECT 99.130 2804.490 100.310 2805.670 ;
        RECT 100.730 2804.490 101.910 2805.670 ;
        RECT 99.130 2626.090 100.310 2627.270 ;
        RECT 100.730 2626.090 101.910 2627.270 ;
        RECT 99.130 2624.490 100.310 2625.670 ;
        RECT 100.730 2624.490 101.910 2625.670 ;
        RECT 99.130 2446.090 100.310 2447.270 ;
        RECT 100.730 2446.090 101.910 2447.270 ;
        RECT 99.130 2444.490 100.310 2445.670 ;
        RECT 100.730 2444.490 101.910 2445.670 ;
        RECT 99.130 2266.090 100.310 2267.270 ;
        RECT 100.730 2266.090 101.910 2267.270 ;
        RECT 99.130 2264.490 100.310 2265.670 ;
        RECT 100.730 2264.490 101.910 2265.670 ;
        RECT 99.130 2086.090 100.310 2087.270 ;
        RECT 100.730 2086.090 101.910 2087.270 ;
        RECT 99.130 2084.490 100.310 2085.670 ;
        RECT 100.730 2084.490 101.910 2085.670 ;
        RECT 99.130 1906.090 100.310 1907.270 ;
        RECT 100.730 1906.090 101.910 1907.270 ;
        RECT 99.130 1904.490 100.310 1905.670 ;
        RECT 100.730 1904.490 101.910 1905.670 ;
        RECT 99.130 1726.090 100.310 1727.270 ;
        RECT 100.730 1726.090 101.910 1727.270 ;
        RECT 99.130 1724.490 100.310 1725.670 ;
        RECT 100.730 1724.490 101.910 1725.670 ;
        RECT 99.130 1546.090 100.310 1547.270 ;
        RECT 100.730 1546.090 101.910 1547.270 ;
        RECT 99.130 1544.490 100.310 1545.670 ;
        RECT 100.730 1544.490 101.910 1545.670 ;
        RECT 99.130 1366.090 100.310 1367.270 ;
        RECT 100.730 1366.090 101.910 1367.270 ;
        RECT 99.130 1364.490 100.310 1365.670 ;
        RECT 100.730 1364.490 101.910 1365.670 ;
        RECT 99.130 1186.090 100.310 1187.270 ;
        RECT 100.730 1186.090 101.910 1187.270 ;
        RECT 99.130 1184.490 100.310 1185.670 ;
        RECT 100.730 1184.490 101.910 1185.670 ;
        RECT 99.130 1006.090 100.310 1007.270 ;
        RECT 100.730 1006.090 101.910 1007.270 ;
        RECT 99.130 1004.490 100.310 1005.670 ;
        RECT 100.730 1004.490 101.910 1005.670 ;
        RECT 99.130 826.090 100.310 827.270 ;
        RECT 100.730 826.090 101.910 827.270 ;
        RECT 99.130 824.490 100.310 825.670 ;
        RECT 100.730 824.490 101.910 825.670 ;
        RECT 99.130 646.090 100.310 647.270 ;
        RECT 100.730 646.090 101.910 647.270 ;
        RECT 99.130 644.490 100.310 645.670 ;
        RECT 100.730 644.490 101.910 645.670 ;
        RECT 99.130 466.090 100.310 467.270 ;
        RECT 100.730 466.090 101.910 467.270 ;
        RECT 99.130 464.490 100.310 465.670 ;
        RECT 100.730 464.490 101.910 465.670 ;
        RECT 99.130 286.090 100.310 287.270 ;
        RECT 100.730 286.090 101.910 287.270 ;
        RECT 99.130 284.490 100.310 285.670 ;
        RECT 100.730 284.490 101.910 285.670 ;
        RECT 99.130 106.090 100.310 107.270 ;
        RECT 100.730 106.090 101.910 107.270 ;
        RECT 99.130 104.490 100.310 105.670 ;
        RECT 100.730 104.490 101.910 105.670 ;
        RECT 99.130 -22.110 100.310 -20.930 ;
        RECT 100.730 -22.110 101.910 -20.930 ;
        RECT 99.130 -23.710 100.310 -22.530 ;
        RECT 100.730 -23.710 101.910 -22.530 ;
        RECT 279.130 3542.210 280.310 3543.390 ;
        RECT 280.730 3542.210 281.910 3543.390 ;
        RECT 279.130 3540.610 280.310 3541.790 ;
        RECT 280.730 3540.610 281.910 3541.790 ;
        RECT 279.130 3346.090 280.310 3347.270 ;
        RECT 280.730 3346.090 281.910 3347.270 ;
        RECT 279.130 3344.490 280.310 3345.670 ;
        RECT 280.730 3344.490 281.910 3345.670 ;
        RECT 279.130 3166.090 280.310 3167.270 ;
        RECT 280.730 3166.090 281.910 3167.270 ;
        RECT 279.130 3164.490 280.310 3165.670 ;
        RECT 280.730 3164.490 281.910 3165.670 ;
        RECT 279.130 2986.090 280.310 2987.270 ;
        RECT 280.730 2986.090 281.910 2987.270 ;
        RECT 279.130 2984.490 280.310 2985.670 ;
        RECT 280.730 2984.490 281.910 2985.670 ;
        RECT 279.130 2806.090 280.310 2807.270 ;
        RECT 280.730 2806.090 281.910 2807.270 ;
        RECT 279.130 2804.490 280.310 2805.670 ;
        RECT 280.730 2804.490 281.910 2805.670 ;
        RECT 279.130 2626.090 280.310 2627.270 ;
        RECT 280.730 2626.090 281.910 2627.270 ;
        RECT 279.130 2624.490 280.310 2625.670 ;
        RECT 280.730 2624.490 281.910 2625.670 ;
        RECT 279.130 2446.090 280.310 2447.270 ;
        RECT 280.730 2446.090 281.910 2447.270 ;
        RECT 279.130 2444.490 280.310 2445.670 ;
        RECT 280.730 2444.490 281.910 2445.670 ;
        RECT 279.130 2266.090 280.310 2267.270 ;
        RECT 280.730 2266.090 281.910 2267.270 ;
        RECT 279.130 2264.490 280.310 2265.670 ;
        RECT 280.730 2264.490 281.910 2265.670 ;
        RECT 279.130 2086.090 280.310 2087.270 ;
        RECT 280.730 2086.090 281.910 2087.270 ;
        RECT 279.130 2084.490 280.310 2085.670 ;
        RECT 280.730 2084.490 281.910 2085.670 ;
        RECT 279.130 1906.090 280.310 1907.270 ;
        RECT 280.730 1906.090 281.910 1907.270 ;
        RECT 279.130 1904.490 280.310 1905.670 ;
        RECT 280.730 1904.490 281.910 1905.670 ;
        RECT 279.130 1726.090 280.310 1727.270 ;
        RECT 280.730 1726.090 281.910 1727.270 ;
        RECT 279.130 1724.490 280.310 1725.670 ;
        RECT 280.730 1724.490 281.910 1725.670 ;
        RECT 279.130 1546.090 280.310 1547.270 ;
        RECT 280.730 1546.090 281.910 1547.270 ;
        RECT 279.130 1544.490 280.310 1545.670 ;
        RECT 280.730 1544.490 281.910 1545.670 ;
        RECT 279.130 1366.090 280.310 1367.270 ;
        RECT 280.730 1366.090 281.910 1367.270 ;
        RECT 279.130 1364.490 280.310 1365.670 ;
        RECT 280.730 1364.490 281.910 1365.670 ;
        RECT 279.130 1186.090 280.310 1187.270 ;
        RECT 280.730 1186.090 281.910 1187.270 ;
        RECT 279.130 1184.490 280.310 1185.670 ;
        RECT 280.730 1184.490 281.910 1185.670 ;
        RECT 279.130 1006.090 280.310 1007.270 ;
        RECT 280.730 1006.090 281.910 1007.270 ;
        RECT 279.130 1004.490 280.310 1005.670 ;
        RECT 280.730 1004.490 281.910 1005.670 ;
        RECT 279.130 826.090 280.310 827.270 ;
        RECT 280.730 826.090 281.910 827.270 ;
        RECT 279.130 824.490 280.310 825.670 ;
        RECT 280.730 824.490 281.910 825.670 ;
        RECT 459.130 3542.210 460.310 3543.390 ;
        RECT 460.730 3542.210 461.910 3543.390 ;
        RECT 459.130 3540.610 460.310 3541.790 ;
        RECT 460.730 3540.610 461.910 3541.790 ;
        RECT 459.130 3346.090 460.310 3347.270 ;
        RECT 460.730 3346.090 461.910 3347.270 ;
        RECT 459.130 3344.490 460.310 3345.670 ;
        RECT 460.730 3344.490 461.910 3345.670 ;
        RECT 459.130 3166.090 460.310 3167.270 ;
        RECT 460.730 3166.090 461.910 3167.270 ;
        RECT 459.130 3164.490 460.310 3165.670 ;
        RECT 460.730 3164.490 461.910 3165.670 ;
        RECT 459.130 2986.090 460.310 2987.270 ;
        RECT 460.730 2986.090 461.910 2987.270 ;
        RECT 459.130 2984.490 460.310 2985.670 ;
        RECT 460.730 2984.490 461.910 2985.670 ;
        RECT 459.130 2806.090 460.310 2807.270 ;
        RECT 460.730 2806.090 461.910 2807.270 ;
        RECT 459.130 2804.490 460.310 2805.670 ;
        RECT 460.730 2804.490 461.910 2805.670 ;
        RECT 459.130 2626.090 460.310 2627.270 ;
        RECT 460.730 2626.090 461.910 2627.270 ;
        RECT 459.130 2624.490 460.310 2625.670 ;
        RECT 460.730 2624.490 461.910 2625.670 ;
        RECT 459.130 2446.090 460.310 2447.270 ;
        RECT 460.730 2446.090 461.910 2447.270 ;
        RECT 459.130 2444.490 460.310 2445.670 ;
        RECT 460.730 2444.490 461.910 2445.670 ;
        RECT 459.130 2266.090 460.310 2267.270 ;
        RECT 460.730 2266.090 461.910 2267.270 ;
        RECT 459.130 2264.490 460.310 2265.670 ;
        RECT 460.730 2264.490 461.910 2265.670 ;
        RECT 459.130 2086.090 460.310 2087.270 ;
        RECT 460.730 2086.090 461.910 2087.270 ;
        RECT 459.130 2084.490 460.310 2085.670 ;
        RECT 460.730 2084.490 461.910 2085.670 ;
        RECT 459.130 1906.090 460.310 1907.270 ;
        RECT 460.730 1906.090 461.910 1907.270 ;
        RECT 459.130 1904.490 460.310 1905.670 ;
        RECT 460.730 1904.490 461.910 1905.670 ;
        RECT 459.130 1726.090 460.310 1727.270 ;
        RECT 460.730 1726.090 461.910 1727.270 ;
        RECT 459.130 1724.490 460.310 1725.670 ;
        RECT 460.730 1724.490 461.910 1725.670 ;
        RECT 459.130 1546.090 460.310 1547.270 ;
        RECT 460.730 1546.090 461.910 1547.270 ;
        RECT 459.130 1544.490 460.310 1545.670 ;
        RECT 460.730 1544.490 461.910 1545.670 ;
        RECT 459.130 1366.090 460.310 1367.270 ;
        RECT 460.730 1366.090 461.910 1367.270 ;
        RECT 459.130 1364.490 460.310 1365.670 ;
        RECT 460.730 1364.490 461.910 1365.670 ;
        RECT 459.130 1186.090 460.310 1187.270 ;
        RECT 460.730 1186.090 461.910 1187.270 ;
        RECT 459.130 1184.490 460.310 1185.670 ;
        RECT 460.730 1184.490 461.910 1185.670 ;
        RECT 459.130 1006.090 460.310 1007.270 ;
        RECT 460.730 1006.090 461.910 1007.270 ;
        RECT 459.130 1004.490 460.310 1005.670 ;
        RECT 460.730 1004.490 461.910 1005.670 ;
        RECT 459.130 826.090 460.310 827.270 ;
        RECT 460.730 826.090 461.910 827.270 ;
        RECT 459.130 824.490 460.310 825.670 ;
        RECT 460.730 824.490 461.910 825.670 ;
        RECT 639.130 3542.210 640.310 3543.390 ;
        RECT 640.730 3542.210 641.910 3543.390 ;
        RECT 639.130 3540.610 640.310 3541.790 ;
        RECT 640.730 3540.610 641.910 3541.790 ;
        RECT 639.130 3346.090 640.310 3347.270 ;
        RECT 640.730 3346.090 641.910 3347.270 ;
        RECT 639.130 3344.490 640.310 3345.670 ;
        RECT 640.730 3344.490 641.910 3345.670 ;
        RECT 639.130 3166.090 640.310 3167.270 ;
        RECT 640.730 3166.090 641.910 3167.270 ;
        RECT 639.130 3164.490 640.310 3165.670 ;
        RECT 640.730 3164.490 641.910 3165.670 ;
        RECT 639.130 2986.090 640.310 2987.270 ;
        RECT 640.730 2986.090 641.910 2987.270 ;
        RECT 639.130 2984.490 640.310 2985.670 ;
        RECT 640.730 2984.490 641.910 2985.670 ;
        RECT 639.130 2806.090 640.310 2807.270 ;
        RECT 640.730 2806.090 641.910 2807.270 ;
        RECT 639.130 2804.490 640.310 2805.670 ;
        RECT 640.730 2804.490 641.910 2805.670 ;
        RECT 639.130 2626.090 640.310 2627.270 ;
        RECT 640.730 2626.090 641.910 2627.270 ;
        RECT 639.130 2624.490 640.310 2625.670 ;
        RECT 640.730 2624.490 641.910 2625.670 ;
        RECT 639.130 2446.090 640.310 2447.270 ;
        RECT 640.730 2446.090 641.910 2447.270 ;
        RECT 639.130 2444.490 640.310 2445.670 ;
        RECT 640.730 2444.490 641.910 2445.670 ;
        RECT 639.130 2266.090 640.310 2267.270 ;
        RECT 640.730 2266.090 641.910 2267.270 ;
        RECT 639.130 2264.490 640.310 2265.670 ;
        RECT 640.730 2264.490 641.910 2265.670 ;
        RECT 639.130 2086.090 640.310 2087.270 ;
        RECT 640.730 2086.090 641.910 2087.270 ;
        RECT 639.130 2084.490 640.310 2085.670 ;
        RECT 640.730 2084.490 641.910 2085.670 ;
        RECT 639.130 1906.090 640.310 1907.270 ;
        RECT 640.730 1906.090 641.910 1907.270 ;
        RECT 639.130 1904.490 640.310 1905.670 ;
        RECT 640.730 1904.490 641.910 1905.670 ;
        RECT 639.130 1726.090 640.310 1727.270 ;
        RECT 640.730 1726.090 641.910 1727.270 ;
        RECT 639.130 1724.490 640.310 1725.670 ;
        RECT 640.730 1724.490 641.910 1725.670 ;
        RECT 639.130 1546.090 640.310 1547.270 ;
        RECT 640.730 1546.090 641.910 1547.270 ;
        RECT 639.130 1544.490 640.310 1545.670 ;
        RECT 640.730 1544.490 641.910 1545.670 ;
        RECT 639.130 1366.090 640.310 1367.270 ;
        RECT 640.730 1366.090 641.910 1367.270 ;
        RECT 639.130 1364.490 640.310 1365.670 ;
        RECT 640.730 1364.490 641.910 1365.670 ;
        RECT 639.130 1186.090 640.310 1187.270 ;
        RECT 640.730 1186.090 641.910 1187.270 ;
        RECT 639.130 1184.490 640.310 1185.670 ;
        RECT 640.730 1184.490 641.910 1185.670 ;
        RECT 639.130 1006.090 640.310 1007.270 ;
        RECT 640.730 1006.090 641.910 1007.270 ;
        RECT 639.130 1004.490 640.310 1005.670 ;
        RECT 640.730 1004.490 641.910 1005.670 ;
        RECT 639.130 826.090 640.310 827.270 ;
        RECT 640.730 826.090 641.910 827.270 ;
        RECT 639.130 824.490 640.310 825.670 ;
        RECT 640.730 824.490 641.910 825.670 ;
        RECT 819.130 3542.210 820.310 3543.390 ;
        RECT 820.730 3542.210 821.910 3543.390 ;
        RECT 819.130 3540.610 820.310 3541.790 ;
        RECT 820.730 3540.610 821.910 3541.790 ;
        RECT 819.130 3346.090 820.310 3347.270 ;
        RECT 820.730 3346.090 821.910 3347.270 ;
        RECT 819.130 3344.490 820.310 3345.670 ;
        RECT 820.730 3344.490 821.910 3345.670 ;
        RECT 819.130 3166.090 820.310 3167.270 ;
        RECT 820.730 3166.090 821.910 3167.270 ;
        RECT 819.130 3164.490 820.310 3165.670 ;
        RECT 820.730 3164.490 821.910 3165.670 ;
        RECT 819.130 2986.090 820.310 2987.270 ;
        RECT 820.730 2986.090 821.910 2987.270 ;
        RECT 819.130 2984.490 820.310 2985.670 ;
        RECT 820.730 2984.490 821.910 2985.670 ;
        RECT 819.130 2806.090 820.310 2807.270 ;
        RECT 820.730 2806.090 821.910 2807.270 ;
        RECT 819.130 2804.490 820.310 2805.670 ;
        RECT 820.730 2804.490 821.910 2805.670 ;
        RECT 819.130 2626.090 820.310 2627.270 ;
        RECT 820.730 2626.090 821.910 2627.270 ;
        RECT 819.130 2624.490 820.310 2625.670 ;
        RECT 820.730 2624.490 821.910 2625.670 ;
        RECT 819.130 2446.090 820.310 2447.270 ;
        RECT 820.730 2446.090 821.910 2447.270 ;
        RECT 819.130 2444.490 820.310 2445.670 ;
        RECT 820.730 2444.490 821.910 2445.670 ;
        RECT 819.130 2266.090 820.310 2267.270 ;
        RECT 820.730 2266.090 821.910 2267.270 ;
        RECT 819.130 2264.490 820.310 2265.670 ;
        RECT 820.730 2264.490 821.910 2265.670 ;
        RECT 819.130 2086.090 820.310 2087.270 ;
        RECT 820.730 2086.090 821.910 2087.270 ;
        RECT 819.130 2084.490 820.310 2085.670 ;
        RECT 820.730 2084.490 821.910 2085.670 ;
        RECT 819.130 1906.090 820.310 1907.270 ;
        RECT 820.730 1906.090 821.910 1907.270 ;
        RECT 819.130 1904.490 820.310 1905.670 ;
        RECT 820.730 1904.490 821.910 1905.670 ;
        RECT 819.130 1726.090 820.310 1727.270 ;
        RECT 820.730 1726.090 821.910 1727.270 ;
        RECT 819.130 1724.490 820.310 1725.670 ;
        RECT 820.730 1724.490 821.910 1725.670 ;
        RECT 819.130 1546.090 820.310 1547.270 ;
        RECT 820.730 1546.090 821.910 1547.270 ;
        RECT 819.130 1544.490 820.310 1545.670 ;
        RECT 820.730 1544.490 821.910 1545.670 ;
        RECT 819.130 1366.090 820.310 1367.270 ;
        RECT 820.730 1366.090 821.910 1367.270 ;
        RECT 819.130 1364.490 820.310 1365.670 ;
        RECT 820.730 1364.490 821.910 1365.670 ;
        RECT 819.130 1186.090 820.310 1187.270 ;
        RECT 820.730 1186.090 821.910 1187.270 ;
        RECT 819.130 1184.490 820.310 1185.670 ;
        RECT 820.730 1184.490 821.910 1185.670 ;
        RECT 819.130 1006.090 820.310 1007.270 ;
        RECT 820.730 1006.090 821.910 1007.270 ;
        RECT 819.130 1004.490 820.310 1005.670 ;
        RECT 820.730 1004.490 821.910 1005.670 ;
        RECT 819.130 826.090 820.310 827.270 ;
        RECT 820.730 826.090 821.910 827.270 ;
        RECT 819.130 824.490 820.310 825.670 ;
        RECT 820.730 824.490 821.910 825.670 ;
        RECT 279.130 646.090 280.310 647.270 ;
        RECT 280.730 646.090 281.910 647.270 ;
        RECT 279.130 644.490 280.310 645.670 ;
        RECT 280.730 644.490 281.910 645.670 ;
        RECT 819.130 646.090 820.310 647.270 ;
        RECT 820.730 646.090 821.910 647.270 ;
        RECT 819.130 644.490 820.310 645.670 ;
        RECT 820.730 644.490 821.910 645.670 ;
        RECT 279.130 466.090 280.310 467.270 ;
        RECT 280.730 466.090 281.910 467.270 ;
        RECT 279.130 464.490 280.310 465.670 ;
        RECT 280.730 464.490 281.910 465.670 ;
        RECT 279.130 286.090 280.310 287.270 ;
        RECT 280.730 286.090 281.910 287.270 ;
        RECT 279.130 284.490 280.310 285.670 ;
        RECT 280.730 284.490 281.910 285.670 ;
        RECT 279.130 106.090 280.310 107.270 ;
        RECT 280.730 106.090 281.910 107.270 ;
        RECT 279.130 104.490 280.310 105.670 ;
        RECT 280.730 104.490 281.910 105.670 ;
        RECT 279.130 -22.110 280.310 -20.930 ;
        RECT 280.730 -22.110 281.910 -20.930 ;
        RECT 279.130 -23.710 280.310 -22.530 ;
        RECT 280.730 -23.710 281.910 -22.530 ;
        RECT 459.130 466.090 460.310 467.270 ;
        RECT 460.730 466.090 461.910 467.270 ;
        RECT 459.130 464.490 460.310 465.670 ;
        RECT 460.730 464.490 461.910 465.670 ;
        RECT 459.130 286.090 460.310 287.270 ;
        RECT 460.730 286.090 461.910 287.270 ;
        RECT 459.130 284.490 460.310 285.670 ;
        RECT 460.730 284.490 461.910 285.670 ;
        RECT 459.130 106.090 460.310 107.270 ;
        RECT 460.730 106.090 461.910 107.270 ;
        RECT 459.130 104.490 460.310 105.670 ;
        RECT 460.730 104.490 461.910 105.670 ;
        RECT 459.130 -22.110 460.310 -20.930 ;
        RECT 460.730 -22.110 461.910 -20.930 ;
        RECT 459.130 -23.710 460.310 -22.530 ;
        RECT 460.730 -23.710 461.910 -22.530 ;
        RECT 639.130 466.090 640.310 467.270 ;
        RECT 640.730 466.090 641.910 467.270 ;
        RECT 639.130 464.490 640.310 465.670 ;
        RECT 640.730 464.490 641.910 465.670 ;
        RECT 639.130 286.090 640.310 287.270 ;
        RECT 640.730 286.090 641.910 287.270 ;
        RECT 639.130 284.490 640.310 285.670 ;
        RECT 640.730 284.490 641.910 285.670 ;
        RECT 639.130 106.090 640.310 107.270 ;
        RECT 640.730 106.090 641.910 107.270 ;
        RECT 639.130 104.490 640.310 105.670 ;
        RECT 640.730 104.490 641.910 105.670 ;
        RECT 639.130 -22.110 640.310 -20.930 ;
        RECT 640.730 -22.110 641.910 -20.930 ;
        RECT 639.130 -23.710 640.310 -22.530 ;
        RECT 640.730 -23.710 641.910 -22.530 ;
        RECT 819.130 466.090 820.310 467.270 ;
        RECT 820.730 466.090 821.910 467.270 ;
        RECT 819.130 464.490 820.310 465.670 ;
        RECT 820.730 464.490 821.910 465.670 ;
        RECT 819.130 286.090 820.310 287.270 ;
        RECT 820.730 286.090 821.910 287.270 ;
        RECT 819.130 284.490 820.310 285.670 ;
        RECT 820.730 284.490 821.910 285.670 ;
        RECT 819.130 106.090 820.310 107.270 ;
        RECT 820.730 106.090 821.910 107.270 ;
        RECT 819.130 104.490 820.310 105.670 ;
        RECT 820.730 104.490 821.910 105.670 ;
        RECT 819.130 -22.110 820.310 -20.930 ;
        RECT 820.730 -22.110 821.910 -20.930 ;
        RECT 819.130 -23.710 820.310 -22.530 ;
        RECT 820.730 -23.710 821.910 -22.530 ;
        RECT 999.130 3542.210 1000.310 3543.390 ;
        RECT 1000.730 3542.210 1001.910 3543.390 ;
        RECT 999.130 3540.610 1000.310 3541.790 ;
        RECT 1000.730 3540.610 1001.910 3541.790 ;
        RECT 999.130 3346.090 1000.310 3347.270 ;
        RECT 1000.730 3346.090 1001.910 3347.270 ;
        RECT 999.130 3344.490 1000.310 3345.670 ;
        RECT 1000.730 3344.490 1001.910 3345.670 ;
        RECT 999.130 3166.090 1000.310 3167.270 ;
        RECT 1000.730 3166.090 1001.910 3167.270 ;
        RECT 999.130 3164.490 1000.310 3165.670 ;
        RECT 1000.730 3164.490 1001.910 3165.670 ;
        RECT 999.130 2986.090 1000.310 2987.270 ;
        RECT 1000.730 2986.090 1001.910 2987.270 ;
        RECT 999.130 2984.490 1000.310 2985.670 ;
        RECT 1000.730 2984.490 1001.910 2985.670 ;
        RECT 999.130 2806.090 1000.310 2807.270 ;
        RECT 1000.730 2806.090 1001.910 2807.270 ;
        RECT 999.130 2804.490 1000.310 2805.670 ;
        RECT 1000.730 2804.490 1001.910 2805.670 ;
        RECT 999.130 2626.090 1000.310 2627.270 ;
        RECT 1000.730 2626.090 1001.910 2627.270 ;
        RECT 999.130 2624.490 1000.310 2625.670 ;
        RECT 1000.730 2624.490 1001.910 2625.670 ;
        RECT 999.130 2446.090 1000.310 2447.270 ;
        RECT 1000.730 2446.090 1001.910 2447.270 ;
        RECT 999.130 2444.490 1000.310 2445.670 ;
        RECT 1000.730 2444.490 1001.910 2445.670 ;
        RECT 999.130 2266.090 1000.310 2267.270 ;
        RECT 1000.730 2266.090 1001.910 2267.270 ;
        RECT 999.130 2264.490 1000.310 2265.670 ;
        RECT 1000.730 2264.490 1001.910 2265.670 ;
        RECT 999.130 2086.090 1000.310 2087.270 ;
        RECT 1000.730 2086.090 1001.910 2087.270 ;
        RECT 999.130 2084.490 1000.310 2085.670 ;
        RECT 1000.730 2084.490 1001.910 2085.670 ;
        RECT 999.130 1906.090 1000.310 1907.270 ;
        RECT 1000.730 1906.090 1001.910 1907.270 ;
        RECT 999.130 1904.490 1000.310 1905.670 ;
        RECT 1000.730 1904.490 1001.910 1905.670 ;
        RECT 999.130 1726.090 1000.310 1727.270 ;
        RECT 1000.730 1726.090 1001.910 1727.270 ;
        RECT 999.130 1724.490 1000.310 1725.670 ;
        RECT 1000.730 1724.490 1001.910 1725.670 ;
        RECT 999.130 1546.090 1000.310 1547.270 ;
        RECT 1000.730 1546.090 1001.910 1547.270 ;
        RECT 999.130 1544.490 1000.310 1545.670 ;
        RECT 1000.730 1544.490 1001.910 1545.670 ;
        RECT 999.130 1366.090 1000.310 1367.270 ;
        RECT 1000.730 1366.090 1001.910 1367.270 ;
        RECT 999.130 1364.490 1000.310 1365.670 ;
        RECT 1000.730 1364.490 1001.910 1365.670 ;
        RECT 999.130 1186.090 1000.310 1187.270 ;
        RECT 1000.730 1186.090 1001.910 1187.270 ;
        RECT 999.130 1184.490 1000.310 1185.670 ;
        RECT 1000.730 1184.490 1001.910 1185.670 ;
        RECT 999.130 1006.090 1000.310 1007.270 ;
        RECT 1000.730 1006.090 1001.910 1007.270 ;
        RECT 999.130 1004.490 1000.310 1005.670 ;
        RECT 1000.730 1004.490 1001.910 1005.670 ;
        RECT 999.130 826.090 1000.310 827.270 ;
        RECT 1000.730 826.090 1001.910 827.270 ;
        RECT 999.130 824.490 1000.310 825.670 ;
        RECT 1000.730 824.490 1001.910 825.670 ;
        RECT 999.130 646.090 1000.310 647.270 ;
        RECT 1000.730 646.090 1001.910 647.270 ;
        RECT 999.130 644.490 1000.310 645.670 ;
        RECT 1000.730 644.490 1001.910 645.670 ;
        RECT 999.130 466.090 1000.310 467.270 ;
        RECT 1000.730 466.090 1001.910 467.270 ;
        RECT 999.130 464.490 1000.310 465.670 ;
        RECT 1000.730 464.490 1001.910 465.670 ;
        RECT 999.130 286.090 1000.310 287.270 ;
        RECT 1000.730 286.090 1001.910 287.270 ;
        RECT 999.130 284.490 1000.310 285.670 ;
        RECT 1000.730 284.490 1001.910 285.670 ;
        RECT 999.130 106.090 1000.310 107.270 ;
        RECT 1000.730 106.090 1001.910 107.270 ;
        RECT 999.130 104.490 1000.310 105.670 ;
        RECT 1000.730 104.490 1001.910 105.670 ;
        RECT 999.130 -22.110 1000.310 -20.930 ;
        RECT 1000.730 -22.110 1001.910 -20.930 ;
        RECT 999.130 -23.710 1000.310 -22.530 ;
        RECT 1000.730 -23.710 1001.910 -22.530 ;
        RECT 1179.130 3542.210 1180.310 3543.390 ;
        RECT 1180.730 3542.210 1181.910 3543.390 ;
        RECT 1179.130 3540.610 1180.310 3541.790 ;
        RECT 1180.730 3540.610 1181.910 3541.790 ;
        RECT 1179.130 3346.090 1180.310 3347.270 ;
        RECT 1180.730 3346.090 1181.910 3347.270 ;
        RECT 1179.130 3344.490 1180.310 3345.670 ;
        RECT 1180.730 3344.490 1181.910 3345.670 ;
        RECT 1179.130 3166.090 1180.310 3167.270 ;
        RECT 1180.730 3166.090 1181.910 3167.270 ;
        RECT 1179.130 3164.490 1180.310 3165.670 ;
        RECT 1180.730 3164.490 1181.910 3165.670 ;
        RECT 1179.130 2986.090 1180.310 2987.270 ;
        RECT 1180.730 2986.090 1181.910 2987.270 ;
        RECT 1179.130 2984.490 1180.310 2985.670 ;
        RECT 1180.730 2984.490 1181.910 2985.670 ;
        RECT 1179.130 2806.090 1180.310 2807.270 ;
        RECT 1180.730 2806.090 1181.910 2807.270 ;
        RECT 1179.130 2804.490 1180.310 2805.670 ;
        RECT 1180.730 2804.490 1181.910 2805.670 ;
        RECT 1179.130 2626.090 1180.310 2627.270 ;
        RECT 1180.730 2626.090 1181.910 2627.270 ;
        RECT 1179.130 2624.490 1180.310 2625.670 ;
        RECT 1180.730 2624.490 1181.910 2625.670 ;
        RECT 1179.130 2446.090 1180.310 2447.270 ;
        RECT 1180.730 2446.090 1181.910 2447.270 ;
        RECT 1179.130 2444.490 1180.310 2445.670 ;
        RECT 1180.730 2444.490 1181.910 2445.670 ;
        RECT 1179.130 2266.090 1180.310 2267.270 ;
        RECT 1180.730 2266.090 1181.910 2267.270 ;
        RECT 1179.130 2264.490 1180.310 2265.670 ;
        RECT 1180.730 2264.490 1181.910 2265.670 ;
        RECT 1179.130 2086.090 1180.310 2087.270 ;
        RECT 1180.730 2086.090 1181.910 2087.270 ;
        RECT 1179.130 2084.490 1180.310 2085.670 ;
        RECT 1180.730 2084.490 1181.910 2085.670 ;
        RECT 1179.130 1906.090 1180.310 1907.270 ;
        RECT 1180.730 1906.090 1181.910 1907.270 ;
        RECT 1179.130 1904.490 1180.310 1905.670 ;
        RECT 1180.730 1904.490 1181.910 1905.670 ;
        RECT 1179.130 1726.090 1180.310 1727.270 ;
        RECT 1180.730 1726.090 1181.910 1727.270 ;
        RECT 1179.130 1724.490 1180.310 1725.670 ;
        RECT 1180.730 1724.490 1181.910 1725.670 ;
        RECT 1179.130 1546.090 1180.310 1547.270 ;
        RECT 1180.730 1546.090 1181.910 1547.270 ;
        RECT 1179.130 1544.490 1180.310 1545.670 ;
        RECT 1180.730 1544.490 1181.910 1545.670 ;
        RECT 1179.130 1366.090 1180.310 1367.270 ;
        RECT 1180.730 1366.090 1181.910 1367.270 ;
        RECT 1179.130 1364.490 1180.310 1365.670 ;
        RECT 1180.730 1364.490 1181.910 1365.670 ;
        RECT 1179.130 1186.090 1180.310 1187.270 ;
        RECT 1180.730 1186.090 1181.910 1187.270 ;
        RECT 1179.130 1184.490 1180.310 1185.670 ;
        RECT 1180.730 1184.490 1181.910 1185.670 ;
        RECT 1179.130 1006.090 1180.310 1007.270 ;
        RECT 1180.730 1006.090 1181.910 1007.270 ;
        RECT 1179.130 1004.490 1180.310 1005.670 ;
        RECT 1180.730 1004.490 1181.910 1005.670 ;
        RECT 1179.130 826.090 1180.310 827.270 ;
        RECT 1180.730 826.090 1181.910 827.270 ;
        RECT 1179.130 824.490 1180.310 825.670 ;
        RECT 1180.730 824.490 1181.910 825.670 ;
        RECT 1179.130 646.090 1180.310 647.270 ;
        RECT 1180.730 646.090 1181.910 647.270 ;
        RECT 1179.130 644.490 1180.310 645.670 ;
        RECT 1180.730 644.490 1181.910 645.670 ;
        RECT 1179.130 466.090 1180.310 467.270 ;
        RECT 1180.730 466.090 1181.910 467.270 ;
        RECT 1179.130 464.490 1180.310 465.670 ;
        RECT 1180.730 464.490 1181.910 465.670 ;
        RECT 1179.130 286.090 1180.310 287.270 ;
        RECT 1180.730 286.090 1181.910 287.270 ;
        RECT 1179.130 284.490 1180.310 285.670 ;
        RECT 1180.730 284.490 1181.910 285.670 ;
        RECT 1179.130 106.090 1180.310 107.270 ;
        RECT 1180.730 106.090 1181.910 107.270 ;
        RECT 1179.130 104.490 1180.310 105.670 ;
        RECT 1180.730 104.490 1181.910 105.670 ;
        RECT 1179.130 -22.110 1180.310 -20.930 ;
        RECT 1180.730 -22.110 1181.910 -20.930 ;
        RECT 1179.130 -23.710 1180.310 -22.530 ;
        RECT 1180.730 -23.710 1181.910 -22.530 ;
        RECT 1359.130 3542.210 1360.310 3543.390 ;
        RECT 1360.730 3542.210 1361.910 3543.390 ;
        RECT 1359.130 3540.610 1360.310 3541.790 ;
        RECT 1360.730 3540.610 1361.910 3541.790 ;
        RECT 1359.130 3346.090 1360.310 3347.270 ;
        RECT 1360.730 3346.090 1361.910 3347.270 ;
        RECT 1359.130 3344.490 1360.310 3345.670 ;
        RECT 1360.730 3344.490 1361.910 3345.670 ;
        RECT 1359.130 3166.090 1360.310 3167.270 ;
        RECT 1360.730 3166.090 1361.910 3167.270 ;
        RECT 1359.130 3164.490 1360.310 3165.670 ;
        RECT 1360.730 3164.490 1361.910 3165.670 ;
        RECT 1359.130 2986.090 1360.310 2987.270 ;
        RECT 1360.730 2986.090 1361.910 2987.270 ;
        RECT 1359.130 2984.490 1360.310 2985.670 ;
        RECT 1360.730 2984.490 1361.910 2985.670 ;
        RECT 1359.130 2806.090 1360.310 2807.270 ;
        RECT 1360.730 2806.090 1361.910 2807.270 ;
        RECT 1359.130 2804.490 1360.310 2805.670 ;
        RECT 1360.730 2804.490 1361.910 2805.670 ;
        RECT 1359.130 2626.090 1360.310 2627.270 ;
        RECT 1360.730 2626.090 1361.910 2627.270 ;
        RECT 1359.130 2624.490 1360.310 2625.670 ;
        RECT 1360.730 2624.490 1361.910 2625.670 ;
        RECT 1359.130 2446.090 1360.310 2447.270 ;
        RECT 1360.730 2446.090 1361.910 2447.270 ;
        RECT 1359.130 2444.490 1360.310 2445.670 ;
        RECT 1360.730 2444.490 1361.910 2445.670 ;
        RECT 1359.130 2266.090 1360.310 2267.270 ;
        RECT 1360.730 2266.090 1361.910 2267.270 ;
        RECT 1359.130 2264.490 1360.310 2265.670 ;
        RECT 1360.730 2264.490 1361.910 2265.670 ;
        RECT 1359.130 2086.090 1360.310 2087.270 ;
        RECT 1360.730 2086.090 1361.910 2087.270 ;
        RECT 1359.130 2084.490 1360.310 2085.670 ;
        RECT 1360.730 2084.490 1361.910 2085.670 ;
        RECT 1359.130 1906.090 1360.310 1907.270 ;
        RECT 1360.730 1906.090 1361.910 1907.270 ;
        RECT 1359.130 1904.490 1360.310 1905.670 ;
        RECT 1360.730 1904.490 1361.910 1905.670 ;
        RECT 1359.130 1726.090 1360.310 1727.270 ;
        RECT 1360.730 1726.090 1361.910 1727.270 ;
        RECT 1359.130 1724.490 1360.310 1725.670 ;
        RECT 1360.730 1724.490 1361.910 1725.670 ;
        RECT 1359.130 1546.090 1360.310 1547.270 ;
        RECT 1360.730 1546.090 1361.910 1547.270 ;
        RECT 1359.130 1544.490 1360.310 1545.670 ;
        RECT 1360.730 1544.490 1361.910 1545.670 ;
        RECT 1359.130 1366.090 1360.310 1367.270 ;
        RECT 1360.730 1366.090 1361.910 1367.270 ;
        RECT 1359.130 1364.490 1360.310 1365.670 ;
        RECT 1360.730 1364.490 1361.910 1365.670 ;
        RECT 1359.130 1186.090 1360.310 1187.270 ;
        RECT 1360.730 1186.090 1361.910 1187.270 ;
        RECT 1359.130 1184.490 1360.310 1185.670 ;
        RECT 1360.730 1184.490 1361.910 1185.670 ;
        RECT 1359.130 1006.090 1360.310 1007.270 ;
        RECT 1360.730 1006.090 1361.910 1007.270 ;
        RECT 1359.130 1004.490 1360.310 1005.670 ;
        RECT 1360.730 1004.490 1361.910 1005.670 ;
        RECT 1359.130 826.090 1360.310 827.270 ;
        RECT 1360.730 826.090 1361.910 827.270 ;
        RECT 1359.130 824.490 1360.310 825.670 ;
        RECT 1360.730 824.490 1361.910 825.670 ;
        RECT 1359.130 646.090 1360.310 647.270 ;
        RECT 1360.730 646.090 1361.910 647.270 ;
        RECT 1359.130 644.490 1360.310 645.670 ;
        RECT 1360.730 644.490 1361.910 645.670 ;
        RECT 1359.130 466.090 1360.310 467.270 ;
        RECT 1360.730 466.090 1361.910 467.270 ;
        RECT 1359.130 464.490 1360.310 465.670 ;
        RECT 1360.730 464.490 1361.910 465.670 ;
        RECT 1359.130 286.090 1360.310 287.270 ;
        RECT 1360.730 286.090 1361.910 287.270 ;
        RECT 1359.130 284.490 1360.310 285.670 ;
        RECT 1360.730 284.490 1361.910 285.670 ;
        RECT 1359.130 106.090 1360.310 107.270 ;
        RECT 1360.730 106.090 1361.910 107.270 ;
        RECT 1359.130 104.490 1360.310 105.670 ;
        RECT 1360.730 104.490 1361.910 105.670 ;
        RECT 1359.130 -22.110 1360.310 -20.930 ;
        RECT 1360.730 -22.110 1361.910 -20.930 ;
        RECT 1359.130 -23.710 1360.310 -22.530 ;
        RECT 1360.730 -23.710 1361.910 -22.530 ;
        RECT 1539.130 3542.210 1540.310 3543.390 ;
        RECT 1540.730 3542.210 1541.910 3543.390 ;
        RECT 1539.130 3540.610 1540.310 3541.790 ;
        RECT 1540.730 3540.610 1541.910 3541.790 ;
        RECT 1539.130 3346.090 1540.310 3347.270 ;
        RECT 1540.730 3346.090 1541.910 3347.270 ;
        RECT 1539.130 3344.490 1540.310 3345.670 ;
        RECT 1540.730 3344.490 1541.910 3345.670 ;
        RECT 1539.130 3166.090 1540.310 3167.270 ;
        RECT 1540.730 3166.090 1541.910 3167.270 ;
        RECT 1539.130 3164.490 1540.310 3165.670 ;
        RECT 1540.730 3164.490 1541.910 3165.670 ;
        RECT 1539.130 2986.090 1540.310 2987.270 ;
        RECT 1540.730 2986.090 1541.910 2987.270 ;
        RECT 1539.130 2984.490 1540.310 2985.670 ;
        RECT 1540.730 2984.490 1541.910 2985.670 ;
        RECT 1539.130 2806.090 1540.310 2807.270 ;
        RECT 1540.730 2806.090 1541.910 2807.270 ;
        RECT 1539.130 2804.490 1540.310 2805.670 ;
        RECT 1540.730 2804.490 1541.910 2805.670 ;
        RECT 1539.130 2626.090 1540.310 2627.270 ;
        RECT 1540.730 2626.090 1541.910 2627.270 ;
        RECT 1539.130 2624.490 1540.310 2625.670 ;
        RECT 1540.730 2624.490 1541.910 2625.670 ;
        RECT 1539.130 2446.090 1540.310 2447.270 ;
        RECT 1540.730 2446.090 1541.910 2447.270 ;
        RECT 1539.130 2444.490 1540.310 2445.670 ;
        RECT 1540.730 2444.490 1541.910 2445.670 ;
        RECT 1539.130 2266.090 1540.310 2267.270 ;
        RECT 1540.730 2266.090 1541.910 2267.270 ;
        RECT 1539.130 2264.490 1540.310 2265.670 ;
        RECT 1540.730 2264.490 1541.910 2265.670 ;
        RECT 1539.130 2086.090 1540.310 2087.270 ;
        RECT 1540.730 2086.090 1541.910 2087.270 ;
        RECT 1539.130 2084.490 1540.310 2085.670 ;
        RECT 1540.730 2084.490 1541.910 2085.670 ;
        RECT 1539.130 1906.090 1540.310 1907.270 ;
        RECT 1540.730 1906.090 1541.910 1907.270 ;
        RECT 1539.130 1904.490 1540.310 1905.670 ;
        RECT 1540.730 1904.490 1541.910 1905.670 ;
        RECT 1539.130 1726.090 1540.310 1727.270 ;
        RECT 1540.730 1726.090 1541.910 1727.270 ;
        RECT 1539.130 1724.490 1540.310 1725.670 ;
        RECT 1540.730 1724.490 1541.910 1725.670 ;
        RECT 1539.130 1546.090 1540.310 1547.270 ;
        RECT 1540.730 1546.090 1541.910 1547.270 ;
        RECT 1539.130 1544.490 1540.310 1545.670 ;
        RECT 1540.730 1544.490 1541.910 1545.670 ;
        RECT 1539.130 1366.090 1540.310 1367.270 ;
        RECT 1540.730 1366.090 1541.910 1367.270 ;
        RECT 1539.130 1364.490 1540.310 1365.670 ;
        RECT 1540.730 1364.490 1541.910 1365.670 ;
        RECT 1539.130 1186.090 1540.310 1187.270 ;
        RECT 1540.730 1186.090 1541.910 1187.270 ;
        RECT 1539.130 1184.490 1540.310 1185.670 ;
        RECT 1540.730 1184.490 1541.910 1185.670 ;
        RECT 1539.130 1006.090 1540.310 1007.270 ;
        RECT 1540.730 1006.090 1541.910 1007.270 ;
        RECT 1539.130 1004.490 1540.310 1005.670 ;
        RECT 1540.730 1004.490 1541.910 1005.670 ;
        RECT 1539.130 826.090 1540.310 827.270 ;
        RECT 1540.730 826.090 1541.910 827.270 ;
        RECT 1539.130 824.490 1540.310 825.670 ;
        RECT 1540.730 824.490 1541.910 825.670 ;
        RECT 1539.130 646.090 1540.310 647.270 ;
        RECT 1540.730 646.090 1541.910 647.270 ;
        RECT 1539.130 644.490 1540.310 645.670 ;
        RECT 1540.730 644.490 1541.910 645.670 ;
        RECT 1539.130 466.090 1540.310 467.270 ;
        RECT 1540.730 466.090 1541.910 467.270 ;
        RECT 1539.130 464.490 1540.310 465.670 ;
        RECT 1540.730 464.490 1541.910 465.670 ;
        RECT 1539.130 286.090 1540.310 287.270 ;
        RECT 1540.730 286.090 1541.910 287.270 ;
        RECT 1539.130 284.490 1540.310 285.670 ;
        RECT 1540.730 284.490 1541.910 285.670 ;
        RECT 1539.130 106.090 1540.310 107.270 ;
        RECT 1540.730 106.090 1541.910 107.270 ;
        RECT 1539.130 104.490 1540.310 105.670 ;
        RECT 1540.730 104.490 1541.910 105.670 ;
        RECT 1539.130 -22.110 1540.310 -20.930 ;
        RECT 1540.730 -22.110 1541.910 -20.930 ;
        RECT 1539.130 -23.710 1540.310 -22.530 ;
        RECT 1540.730 -23.710 1541.910 -22.530 ;
        RECT 1719.130 3542.210 1720.310 3543.390 ;
        RECT 1720.730 3542.210 1721.910 3543.390 ;
        RECT 1719.130 3540.610 1720.310 3541.790 ;
        RECT 1720.730 3540.610 1721.910 3541.790 ;
        RECT 1719.130 3346.090 1720.310 3347.270 ;
        RECT 1720.730 3346.090 1721.910 3347.270 ;
        RECT 1719.130 3344.490 1720.310 3345.670 ;
        RECT 1720.730 3344.490 1721.910 3345.670 ;
        RECT 1719.130 3166.090 1720.310 3167.270 ;
        RECT 1720.730 3166.090 1721.910 3167.270 ;
        RECT 1719.130 3164.490 1720.310 3165.670 ;
        RECT 1720.730 3164.490 1721.910 3165.670 ;
        RECT 1719.130 2986.090 1720.310 2987.270 ;
        RECT 1720.730 2986.090 1721.910 2987.270 ;
        RECT 1719.130 2984.490 1720.310 2985.670 ;
        RECT 1720.730 2984.490 1721.910 2985.670 ;
        RECT 1719.130 2806.090 1720.310 2807.270 ;
        RECT 1720.730 2806.090 1721.910 2807.270 ;
        RECT 1719.130 2804.490 1720.310 2805.670 ;
        RECT 1720.730 2804.490 1721.910 2805.670 ;
        RECT 1719.130 2626.090 1720.310 2627.270 ;
        RECT 1720.730 2626.090 1721.910 2627.270 ;
        RECT 1719.130 2624.490 1720.310 2625.670 ;
        RECT 1720.730 2624.490 1721.910 2625.670 ;
        RECT 1719.130 2446.090 1720.310 2447.270 ;
        RECT 1720.730 2446.090 1721.910 2447.270 ;
        RECT 1719.130 2444.490 1720.310 2445.670 ;
        RECT 1720.730 2444.490 1721.910 2445.670 ;
        RECT 1719.130 2266.090 1720.310 2267.270 ;
        RECT 1720.730 2266.090 1721.910 2267.270 ;
        RECT 1719.130 2264.490 1720.310 2265.670 ;
        RECT 1720.730 2264.490 1721.910 2265.670 ;
        RECT 1719.130 2086.090 1720.310 2087.270 ;
        RECT 1720.730 2086.090 1721.910 2087.270 ;
        RECT 1719.130 2084.490 1720.310 2085.670 ;
        RECT 1720.730 2084.490 1721.910 2085.670 ;
        RECT 1719.130 1906.090 1720.310 1907.270 ;
        RECT 1720.730 1906.090 1721.910 1907.270 ;
        RECT 1719.130 1904.490 1720.310 1905.670 ;
        RECT 1720.730 1904.490 1721.910 1905.670 ;
        RECT 1719.130 1726.090 1720.310 1727.270 ;
        RECT 1720.730 1726.090 1721.910 1727.270 ;
        RECT 1719.130 1724.490 1720.310 1725.670 ;
        RECT 1720.730 1724.490 1721.910 1725.670 ;
        RECT 1719.130 1546.090 1720.310 1547.270 ;
        RECT 1720.730 1546.090 1721.910 1547.270 ;
        RECT 1719.130 1544.490 1720.310 1545.670 ;
        RECT 1720.730 1544.490 1721.910 1545.670 ;
        RECT 1719.130 1366.090 1720.310 1367.270 ;
        RECT 1720.730 1366.090 1721.910 1367.270 ;
        RECT 1719.130 1364.490 1720.310 1365.670 ;
        RECT 1720.730 1364.490 1721.910 1365.670 ;
        RECT 1719.130 1186.090 1720.310 1187.270 ;
        RECT 1720.730 1186.090 1721.910 1187.270 ;
        RECT 1719.130 1184.490 1720.310 1185.670 ;
        RECT 1720.730 1184.490 1721.910 1185.670 ;
        RECT 1719.130 1006.090 1720.310 1007.270 ;
        RECT 1720.730 1006.090 1721.910 1007.270 ;
        RECT 1719.130 1004.490 1720.310 1005.670 ;
        RECT 1720.730 1004.490 1721.910 1005.670 ;
        RECT 1719.130 826.090 1720.310 827.270 ;
        RECT 1720.730 826.090 1721.910 827.270 ;
        RECT 1719.130 824.490 1720.310 825.670 ;
        RECT 1720.730 824.490 1721.910 825.670 ;
        RECT 1719.130 646.090 1720.310 647.270 ;
        RECT 1720.730 646.090 1721.910 647.270 ;
        RECT 1719.130 644.490 1720.310 645.670 ;
        RECT 1720.730 644.490 1721.910 645.670 ;
        RECT 1719.130 466.090 1720.310 467.270 ;
        RECT 1720.730 466.090 1721.910 467.270 ;
        RECT 1719.130 464.490 1720.310 465.670 ;
        RECT 1720.730 464.490 1721.910 465.670 ;
        RECT 1719.130 286.090 1720.310 287.270 ;
        RECT 1720.730 286.090 1721.910 287.270 ;
        RECT 1719.130 284.490 1720.310 285.670 ;
        RECT 1720.730 284.490 1721.910 285.670 ;
        RECT 1719.130 106.090 1720.310 107.270 ;
        RECT 1720.730 106.090 1721.910 107.270 ;
        RECT 1719.130 104.490 1720.310 105.670 ;
        RECT 1720.730 104.490 1721.910 105.670 ;
        RECT 1719.130 -22.110 1720.310 -20.930 ;
        RECT 1720.730 -22.110 1721.910 -20.930 ;
        RECT 1719.130 -23.710 1720.310 -22.530 ;
        RECT 1720.730 -23.710 1721.910 -22.530 ;
        RECT 1899.130 3542.210 1900.310 3543.390 ;
        RECT 1900.730 3542.210 1901.910 3543.390 ;
        RECT 1899.130 3540.610 1900.310 3541.790 ;
        RECT 1900.730 3540.610 1901.910 3541.790 ;
        RECT 1899.130 3346.090 1900.310 3347.270 ;
        RECT 1900.730 3346.090 1901.910 3347.270 ;
        RECT 1899.130 3344.490 1900.310 3345.670 ;
        RECT 1900.730 3344.490 1901.910 3345.670 ;
        RECT 1899.130 3166.090 1900.310 3167.270 ;
        RECT 1900.730 3166.090 1901.910 3167.270 ;
        RECT 1899.130 3164.490 1900.310 3165.670 ;
        RECT 1900.730 3164.490 1901.910 3165.670 ;
        RECT 1899.130 2986.090 1900.310 2987.270 ;
        RECT 1900.730 2986.090 1901.910 2987.270 ;
        RECT 1899.130 2984.490 1900.310 2985.670 ;
        RECT 1900.730 2984.490 1901.910 2985.670 ;
        RECT 1899.130 2806.090 1900.310 2807.270 ;
        RECT 1900.730 2806.090 1901.910 2807.270 ;
        RECT 1899.130 2804.490 1900.310 2805.670 ;
        RECT 1900.730 2804.490 1901.910 2805.670 ;
        RECT 1899.130 2626.090 1900.310 2627.270 ;
        RECT 1900.730 2626.090 1901.910 2627.270 ;
        RECT 1899.130 2624.490 1900.310 2625.670 ;
        RECT 1900.730 2624.490 1901.910 2625.670 ;
        RECT 1899.130 2446.090 1900.310 2447.270 ;
        RECT 1900.730 2446.090 1901.910 2447.270 ;
        RECT 1899.130 2444.490 1900.310 2445.670 ;
        RECT 1900.730 2444.490 1901.910 2445.670 ;
        RECT 1899.130 2266.090 1900.310 2267.270 ;
        RECT 1900.730 2266.090 1901.910 2267.270 ;
        RECT 1899.130 2264.490 1900.310 2265.670 ;
        RECT 1900.730 2264.490 1901.910 2265.670 ;
        RECT 1899.130 2086.090 1900.310 2087.270 ;
        RECT 1900.730 2086.090 1901.910 2087.270 ;
        RECT 1899.130 2084.490 1900.310 2085.670 ;
        RECT 1900.730 2084.490 1901.910 2085.670 ;
        RECT 1899.130 1906.090 1900.310 1907.270 ;
        RECT 1900.730 1906.090 1901.910 1907.270 ;
        RECT 1899.130 1904.490 1900.310 1905.670 ;
        RECT 1900.730 1904.490 1901.910 1905.670 ;
        RECT 1899.130 1726.090 1900.310 1727.270 ;
        RECT 1900.730 1726.090 1901.910 1727.270 ;
        RECT 1899.130 1724.490 1900.310 1725.670 ;
        RECT 1900.730 1724.490 1901.910 1725.670 ;
        RECT 1899.130 1546.090 1900.310 1547.270 ;
        RECT 1900.730 1546.090 1901.910 1547.270 ;
        RECT 1899.130 1544.490 1900.310 1545.670 ;
        RECT 1900.730 1544.490 1901.910 1545.670 ;
        RECT 1899.130 1366.090 1900.310 1367.270 ;
        RECT 1900.730 1366.090 1901.910 1367.270 ;
        RECT 1899.130 1364.490 1900.310 1365.670 ;
        RECT 1900.730 1364.490 1901.910 1365.670 ;
        RECT 1899.130 1186.090 1900.310 1187.270 ;
        RECT 1900.730 1186.090 1901.910 1187.270 ;
        RECT 1899.130 1184.490 1900.310 1185.670 ;
        RECT 1900.730 1184.490 1901.910 1185.670 ;
        RECT 1899.130 1006.090 1900.310 1007.270 ;
        RECT 1900.730 1006.090 1901.910 1007.270 ;
        RECT 1899.130 1004.490 1900.310 1005.670 ;
        RECT 1900.730 1004.490 1901.910 1005.670 ;
        RECT 1899.130 826.090 1900.310 827.270 ;
        RECT 1900.730 826.090 1901.910 827.270 ;
        RECT 1899.130 824.490 1900.310 825.670 ;
        RECT 1900.730 824.490 1901.910 825.670 ;
        RECT 1899.130 646.090 1900.310 647.270 ;
        RECT 1900.730 646.090 1901.910 647.270 ;
        RECT 1899.130 644.490 1900.310 645.670 ;
        RECT 1900.730 644.490 1901.910 645.670 ;
        RECT 1899.130 466.090 1900.310 467.270 ;
        RECT 1900.730 466.090 1901.910 467.270 ;
        RECT 1899.130 464.490 1900.310 465.670 ;
        RECT 1900.730 464.490 1901.910 465.670 ;
        RECT 1899.130 286.090 1900.310 287.270 ;
        RECT 1900.730 286.090 1901.910 287.270 ;
        RECT 1899.130 284.490 1900.310 285.670 ;
        RECT 1900.730 284.490 1901.910 285.670 ;
        RECT 1899.130 106.090 1900.310 107.270 ;
        RECT 1900.730 106.090 1901.910 107.270 ;
        RECT 1899.130 104.490 1900.310 105.670 ;
        RECT 1900.730 104.490 1901.910 105.670 ;
        RECT 1899.130 -22.110 1900.310 -20.930 ;
        RECT 1900.730 -22.110 1901.910 -20.930 ;
        RECT 1899.130 -23.710 1900.310 -22.530 ;
        RECT 1900.730 -23.710 1901.910 -22.530 ;
        RECT 2079.130 3542.210 2080.310 3543.390 ;
        RECT 2080.730 3542.210 2081.910 3543.390 ;
        RECT 2079.130 3540.610 2080.310 3541.790 ;
        RECT 2080.730 3540.610 2081.910 3541.790 ;
        RECT 2079.130 3346.090 2080.310 3347.270 ;
        RECT 2080.730 3346.090 2081.910 3347.270 ;
        RECT 2079.130 3344.490 2080.310 3345.670 ;
        RECT 2080.730 3344.490 2081.910 3345.670 ;
        RECT 2079.130 3166.090 2080.310 3167.270 ;
        RECT 2080.730 3166.090 2081.910 3167.270 ;
        RECT 2079.130 3164.490 2080.310 3165.670 ;
        RECT 2080.730 3164.490 2081.910 3165.670 ;
        RECT 2079.130 2986.090 2080.310 2987.270 ;
        RECT 2080.730 2986.090 2081.910 2987.270 ;
        RECT 2079.130 2984.490 2080.310 2985.670 ;
        RECT 2080.730 2984.490 2081.910 2985.670 ;
        RECT 2079.130 2806.090 2080.310 2807.270 ;
        RECT 2080.730 2806.090 2081.910 2807.270 ;
        RECT 2079.130 2804.490 2080.310 2805.670 ;
        RECT 2080.730 2804.490 2081.910 2805.670 ;
        RECT 2079.130 2626.090 2080.310 2627.270 ;
        RECT 2080.730 2626.090 2081.910 2627.270 ;
        RECT 2079.130 2624.490 2080.310 2625.670 ;
        RECT 2080.730 2624.490 2081.910 2625.670 ;
        RECT 2079.130 2446.090 2080.310 2447.270 ;
        RECT 2080.730 2446.090 2081.910 2447.270 ;
        RECT 2079.130 2444.490 2080.310 2445.670 ;
        RECT 2080.730 2444.490 2081.910 2445.670 ;
        RECT 2079.130 2266.090 2080.310 2267.270 ;
        RECT 2080.730 2266.090 2081.910 2267.270 ;
        RECT 2079.130 2264.490 2080.310 2265.670 ;
        RECT 2080.730 2264.490 2081.910 2265.670 ;
        RECT 2079.130 2086.090 2080.310 2087.270 ;
        RECT 2080.730 2086.090 2081.910 2087.270 ;
        RECT 2079.130 2084.490 2080.310 2085.670 ;
        RECT 2080.730 2084.490 2081.910 2085.670 ;
        RECT 2079.130 1906.090 2080.310 1907.270 ;
        RECT 2080.730 1906.090 2081.910 1907.270 ;
        RECT 2079.130 1904.490 2080.310 1905.670 ;
        RECT 2080.730 1904.490 2081.910 1905.670 ;
        RECT 2079.130 1726.090 2080.310 1727.270 ;
        RECT 2080.730 1726.090 2081.910 1727.270 ;
        RECT 2079.130 1724.490 2080.310 1725.670 ;
        RECT 2080.730 1724.490 2081.910 1725.670 ;
        RECT 2079.130 1546.090 2080.310 1547.270 ;
        RECT 2080.730 1546.090 2081.910 1547.270 ;
        RECT 2079.130 1544.490 2080.310 1545.670 ;
        RECT 2080.730 1544.490 2081.910 1545.670 ;
        RECT 2079.130 1366.090 2080.310 1367.270 ;
        RECT 2080.730 1366.090 2081.910 1367.270 ;
        RECT 2079.130 1364.490 2080.310 1365.670 ;
        RECT 2080.730 1364.490 2081.910 1365.670 ;
        RECT 2079.130 1186.090 2080.310 1187.270 ;
        RECT 2080.730 1186.090 2081.910 1187.270 ;
        RECT 2079.130 1184.490 2080.310 1185.670 ;
        RECT 2080.730 1184.490 2081.910 1185.670 ;
        RECT 2079.130 1006.090 2080.310 1007.270 ;
        RECT 2080.730 1006.090 2081.910 1007.270 ;
        RECT 2079.130 1004.490 2080.310 1005.670 ;
        RECT 2080.730 1004.490 2081.910 1005.670 ;
        RECT 2079.130 826.090 2080.310 827.270 ;
        RECT 2080.730 826.090 2081.910 827.270 ;
        RECT 2079.130 824.490 2080.310 825.670 ;
        RECT 2080.730 824.490 2081.910 825.670 ;
        RECT 2079.130 646.090 2080.310 647.270 ;
        RECT 2080.730 646.090 2081.910 647.270 ;
        RECT 2079.130 644.490 2080.310 645.670 ;
        RECT 2080.730 644.490 2081.910 645.670 ;
        RECT 2079.130 466.090 2080.310 467.270 ;
        RECT 2080.730 466.090 2081.910 467.270 ;
        RECT 2079.130 464.490 2080.310 465.670 ;
        RECT 2080.730 464.490 2081.910 465.670 ;
        RECT 2079.130 286.090 2080.310 287.270 ;
        RECT 2080.730 286.090 2081.910 287.270 ;
        RECT 2079.130 284.490 2080.310 285.670 ;
        RECT 2080.730 284.490 2081.910 285.670 ;
        RECT 2079.130 106.090 2080.310 107.270 ;
        RECT 2080.730 106.090 2081.910 107.270 ;
        RECT 2079.130 104.490 2080.310 105.670 ;
        RECT 2080.730 104.490 2081.910 105.670 ;
        RECT 2079.130 -22.110 2080.310 -20.930 ;
        RECT 2080.730 -22.110 2081.910 -20.930 ;
        RECT 2079.130 -23.710 2080.310 -22.530 ;
        RECT 2080.730 -23.710 2081.910 -22.530 ;
        RECT 2259.130 3542.210 2260.310 3543.390 ;
        RECT 2260.730 3542.210 2261.910 3543.390 ;
        RECT 2259.130 3540.610 2260.310 3541.790 ;
        RECT 2260.730 3540.610 2261.910 3541.790 ;
        RECT 2259.130 3346.090 2260.310 3347.270 ;
        RECT 2260.730 3346.090 2261.910 3347.270 ;
        RECT 2259.130 3344.490 2260.310 3345.670 ;
        RECT 2260.730 3344.490 2261.910 3345.670 ;
        RECT 2259.130 3166.090 2260.310 3167.270 ;
        RECT 2260.730 3166.090 2261.910 3167.270 ;
        RECT 2259.130 3164.490 2260.310 3165.670 ;
        RECT 2260.730 3164.490 2261.910 3165.670 ;
        RECT 2259.130 2986.090 2260.310 2987.270 ;
        RECT 2260.730 2986.090 2261.910 2987.270 ;
        RECT 2259.130 2984.490 2260.310 2985.670 ;
        RECT 2260.730 2984.490 2261.910 2985.670 ;
        RECT 2259.130 2806.090 2260.310 2807.270 ;
        RECT 2260.730 2806.090 2261.910 2807.270 ;
        RECT 2259.130 2804.490 2260.310 2805.670 ;
        RECT 2260.730 2804.490 2261.910 2805.670 ;
        RECT 2259.130 2626.090 2260.310 2627.270 ;
        RECT 2260.730 2626.090 2261.910 2627.270 ;
        RECT 2259.130 2624.490 2260.310 2625.670 ;
        RECT 2260.730 2624.490 2261.910 2625.670 ;
        RECT 2259.130 2446.090 2260.310 2447.270 ;
        RECT 2260.730 2446.090 2261.910 2447.270 ;
        RECT 2259.130 2444.490 2260.310 2445.670 ;
        RECT 2260.730 2444.490 2261.910 2445.670 ;
        RECT 2259.130 2266.090 2260.310 2267.270 ;
        RECT 2260.730 2266.090 2261.910 2267.270 ;
        RECT 2259.130 2264.490 2260.310 2265.670 ;
        RECT 2260.730 2264.490 2261.910 2265.670 ;
        RECT 2259.130 2086.090 2260.310 2087.270 ;
        RECT 2260.730 2086.090 2261.910 2087.270 ;
        RECT 2259.130 2084.490 2260.310 2085.670 ;
        RECT 2260.730 2084.490 2261.910 2085.670 ;
        RECT 2259.130 1906.090 2260.310 1907.270 ;
        RECT 2260.730 1906.090 2261.910 1907.270 ;
        RECT 2259.130 1904.490 2260.310 1905.670 ;
        RECT 2260.730 1904.490 2261.910 1905.670 ;
        RECT 2259.130 1726.090 2260.310 1727.270 ;
        RECT 2260.730 1726.090 2261.910 1727.270 ;
        RECT 2259.130 1724.490 2260.310 1725.670 ;
        RECT 2260.730 1724.490 2261.910 1725.670 ;
        RECT 2259.130 1546.090 2260.310 1547.270 ;
        RECT 2260.730 1546.090 2261.910 1547.270 ;
        RECT 2259.130 1544.490 2260.310 1545.670 ;
        RECT 2260.730 1544.490 2261.910 1545.670 ;
        RECT 2259.130 1366.090 2260.310 1367.270 ;
        RECT 2260.730 1366.090 2261.910 1367.270 ;
        RECT 2259.130 1364.490 2260.310 1365.670 ;
        RECT 2260.730 1364.490 2261.910 1365.670 ;
        RECT 2259.130 1186.090 2260.310 1187.270 ;
        RECT 2260.730 1186.090 2261.910 1187.270 ;
        RECT 2259.130 1184.490 2260.310 1185.670 ;
        RECT 2260.730 1184.490 2261.910 1185.670 ;
        RECT 2259.130 1006.090 2260.310 1007.270 ;
        RECT 2260.730 1006.090 2261.910 1007.270 ;
        RECT 2259.130 1004.490 2260.310 1005.670 ;
        RECT 2260.730 1004.490 2261.910 1005.670 ;
        RECT 2259.130 826.090 2260.310 827.270 ;
        RECT 2260.730 826.090 2261.910 827.270 ;
        RECT 2259.130 824.490 2260.310 825.670 ;
        RECT 2260.730 824.490 2261.910 825.670 ;
        RECT 2259.130 646.090 2260.310 647.270 ;
        RECT 2260.730 646.090 2261.910 647.270 ;
        RECT 2259.130 644.490 2260.310 645.670 ;
        RECT 2260.730 644.490 2261.910 645.670 ;
        RECT 2259.130 466.090 2260.310 467.270 ;
        RECT 2260.730 466.090 2261.910 467.270 ;
        RECT 2259.130 464.490 2260.310 465.670 ;
        RECT 2260.730 464.490 2261.910 465.670 ;
        RECT 2259.130 286.090 2260.310 287.270 ;
        RECT 2260.730 286.090 2261.910 287.270 ;
        RECT 2259.130 284.490 2260.310 285.670 ;
        RECT 2260.730 284.490 2261.910 285.670 ;
        RECT 2259.130 106.090 2260.310 107.270 ;
        RECT 2260.730 106.090 2261.910 107.270 ;
        RECT 2259.130 104.490 2260.310 105.670 ;
        RECT 2260.730 104.490 2261.910 105.670 ;
        RECT 2259.130 -22.110 2260.310 -20.930 ;
        RECT 2260.730 -22.110 2261.910 -20.930 ;
        RECT 2259.130 -23.710 2260.310 -22.530 ;
        RECT 2260.730 -23.710 2261.910 -22.530 ;
        RECT 2439.130 3542.210 2440.310 3543.390 ;
        RECT 2440.730 3542.210 2441.910 3543.390 ;
        RECT 2439.130 3540.610 2440.310 3541.790 ;
        RECT 2440.730 3540.610 2441.910 3541.790 ;
        RECT 2439.130 3346.090 2440.310 3347.270 ;
        RECT 2440.730 3346.090 2441.910 3347.270 ;
        RECT 2439.130 3344.490 2440.310 3345.670 ;
        RECT 2440.730 3344.490 2441.910 3345.670 ;
        RECT 2439.130 3166.090 2440.310 3167.270 ;
        RECT 2440.730 3166.090 2441.910 3167.270 ;
        RECT 2439.130 3164.490 2440.310 3165.670 ;
        RECT 2440.730 3164.490 2441.910 3165.670 ;
        RECT 2439.130 2986.090 2440.310 2987.270 ;
        RECT 2440.730 2986.090 2441.910 2987.270 ;
        RECT 2439.130 2984.490 2440.310 2985.670 ;
        RECT 2440.730 2984.490 2441.910 2985.670 ;
        RECT 2439.130 2806.090 2440.310 2807.270 ;
        RECT 2440.730 2806.090 2441.910 2807.270 ;
        RECT 2439.130 2804.490 2440.310 2805.670 ;
        RECT 2440.730 2804.490 2441.910 2805.670 ;
        RECT 2439.130 2626.090 2440.310 2627.270 ;
        RECT 2440.730 2626.090 2441.910 2627.270 ;
        RECT 2439.130 2624.490 2440.310 2625.670 ;
        RECT 2440.730 2624.490 2441.910 2625.670 ;
        RECT 2439.130 2446.090 2440.310 2447.270 ;
        RECT 2440.730 2446.090 2441.910 2447.270 ;
        RECT 2439.130 2444.490 2440.310 2445.670 ;
        RECT 2440.730 2444.490 2441.910 2445.670 ;
        RECT 2439.130 2266.090 2440.310 2267.270 ;
        RECT 2440.730 2266.090 2441.910 2267.270 ;
        RECT 2439.130 2264.490 2440.310 2265.670 ;
        RECT 2440.730 2264.490 2441.910 2265.670 ;
        RECT 2439.130 2086.090 2440.310 2087.270 ;
        RECT 2440.730 2086.090 2441.910 2087.270 ;
        RECT 2439.130 2084.490 2440.310 2085.670 ;
        RECT 2440.730 2084.490 2441.910 2085.670 ;
        RECT 2439.130 1906.090 2440.310 1907.270 ;
        RECT 2440.730 1906.090 2441.910 1907.270 ;
        RECT 2439.130 1904.490 2440.310 1905.670 ;
        RECT 2440.730 1904.490 2441.910 1905.670 ;
        RECT 2439.130 1726.090 2440.310 1727.270 ;
        RECT 2440.730 1726.090 2441.910 1727.270 ;
        RECT 2439.130 1724.490 2440.310 1725.670 ;
        RECT 2440.730 1724.490 2441.910 1725.670 ;
        RECT 2439.130 1546.090 2440.310 1547.270 ;
        RECT 2440.730 1546.090 2441.910 1547.270 ;
        RECT 2439.130 1544.490 2440.310 1545.670 ;
        RECT 2440.730 1544.490 2441.910 1545.670 ;
        RECT 2439.130 1366.090 2440.310 1367.270 ;
        RECT 2440.730 1366.090 2441.910 1367.270 ;
        RECT 2439.130 1364.490 2440.310 1365.670 ;
        RECT 2440.730 1364.490 2441.910 1365.670 ;
        RECT 2439.130 1186.090 2440.310 1187.270 ;
        RECT 2440.730 1186.090 2441.910 1187.270 ;
        RECT 2439.130 1184.490 2440.310 1185.670 ;
        RECT 2440.730 1184.490 2441.910 1185.670 ;
        RECT 2439.130 1006.090 2440.310 1007.270 ;
        RECT 2440.730 1006.090 2441.910 1007.270 ;
        RECT 2439.130 1004.490 2440.310 1005.670 ;
        RECT 2440.730 1004.490 2441.910 1005.670 ;
        RECT 2439.130 826.090 2440.310 827.270 ;
        RECT 2440.730 826.090 2441.910 827.270 ;
        RECT 2439.130 824.490 2440.310 825.670 ;
        RECT 2440.730 824.490 2441.910 825.670 ;
        RECT 2439.130 646.090 2440.310 647.270 ;
        RECT 2440.730 646.090 2441.910 647.270 ;
        RECT 2439.130 644.490 2440.310 645.670 ;
        RECT 2440.730 644.490 2441.910 645.670 ;
        RECT 2439.130 466.090 2440.310 467.270 ;
        RECT 2440.730 466.090 2441.910 467.270 ;
        RECT 2439.130 464.490 2440.310 465.670 ;
        RECT 2440.730 464.490 2441.910 465.670 ;
        RECT 2439.130 286.090 2440.310 287.270 ;
        RECT 2440.730 286.090 2441.910 287.270 ;
        RECT 2439.130 284.490 2440.310 285.670 ;
        RECT 2440.730 284.490 2441.910 285.670 ;
        RECT 2439.130 106.090 2440.310 107.270 ;
        RECT 2440.730 106.090 2441.910 107.270 ;
        RECT 2439.130 104.490 2440.310 105.670 ;
        RECT 2440.730 104.490 2441.910 105.670 ;
        RECT 2439.130 -22.110 2440.310 -20.930 ;
        RECT 2440.730 -22.110 2441.910 -20.930 ;
        RECT 2439.130 -23.710 2440.310 -22.530 ;
        RECT 2440.730 -23.710 2441.910 -22.530 ;
        RECT 2619.130 3542.210 2620.310 3543.390 ;
        RECT 2620.730 3542.210 2621.910 3543.390 ;
        RECT 2619.130 3540.610 2620.310 3541.790 ;
        RECT 2620.730 3540.610 2621.910 3541.790 ;
        RECT 2619.130 3346.090 2620.310 3347.270 ;
        RECT 2620.730 3346.090 2621.910 3347.270 ;
        RECT 2619.130 3344.490 2620.310 3345.670 ;
        RECT 2620.730 3344.490 2621.910 3345.670 ;
        RECT 2619.130 3166.090 2620.310 3167.270 ;
        RECT 2620.730 3166.090 2621.910 3167.270 ;
        RECT 2619.130 3164.490 2620.310 3165.670 ;
        RECT 2620.730 3164.490 2621.910 3165.670 ;
        RECT 2619.130 2986.090 2620.310 2987.270 ;
        RECT 2620.730 2986.090 2621.910 2987.270 ;
        RECT 2619.130 2984.490 2620.310 2985.670 ;
        RECT 2620.730 2984.490 2621.910 2985.670 ;
        RECT 2619.130 2806.090 2620.310 2807.270 ;
        RECT 2620.730 2806.090 2621.910 2807.270 ;
        RECT 2619.130 2804.490 2620.310 2805.670 ;
        RECT 2620.730 2804.490 2621.910 2805.670 ;
        RECT 2619.130 2626.090 2620.310 2627.270 ;
        RECT 2620.730 2626.090 2621.910 2627.270 ;
        RECT 2619.130 2624.490 2620.310 2625.670 ;
        RECT 2620.730 2624.490 2621.910 2625.670 ;
        RECT 2619.130 2446.090 2620.310 2447.270 ;
        RECT 2620.730 2446.090 2621.910 2447.270 ;
        RECT 2619.130 2444.490 2620.310 2445.670 ;
        RECT 2620.730 2444.490 2621.910 2445.670 ;
        RECT 2619.130 2266.090 2620.310 2267.270 ;
        RECT 2620.730 2266.090 2621.910 2267.270 ;
        RECT 2619.130 2264.490 2620.310 2265.670 ;
        RECT 2620.730 2264.490 2621.910 2265.670 ;
        RECT 2619.130 2086.090 2620.310 2087.270 ;
        RECT 2620.730 2086.090 2621.910 2087.270 ;
        RECT 2619.130 2084.490 2620.310 2085.670 ;
        RECT 2620.730 2084.490 2621.910 2085.670 ;
        RECT 2619.130 1906.090 2620.310 1907.270 ;
        RECT 2620.730 1906.090 2621.910 1907.270 ;
        RECT 2619.130 1904.490 2620.310 1905.670 ;
        RECT 2620.730 1904.490 2621.910 1905.670 ;
        RECT 2619.130 1726.090 2620.310 1727.270 ;
        RECT 2620.730 1726.090 2621.910 1727.270 ;
        RECT 2619.130 1724.490 2620.310 1725.670 ;
        RECT 2620.730 1724.490 2621.910 1725.670 ;
        RECT 2619.130 1546.090 2620.310 1547.270 ;
        RECT 2620.730 1546.090 2621.910 1547.270 ;
        RECT 2619.130 1544.490 2620.310 1545.670 ;
        RECT 2620.730 1544.490 2621.910 1545.670 ;
        RECT 2619.130 1366.090 2620.310 1367.270 ;
        RECT 2620.730 1366.090 2621.910 1367.270 ;
        RECT 2619.130 1364.490 2620.310 1365.670 ;
        RECT 2620.730 1364.490 2621.910 1365.670 ;
        RECT 2619.130 1186.090 2620.310 1187.270 ;
        RECT 2620.730 1186.090 2621.910 1187.270 ;
        RECT 2619.130 1184.490 2620.310 1185.670 ;
        RECT 2620.730 1184.490 2621.910 1185.670 ;
        RECT 2619.130 1006.090 2620.310 1007.270 ;
        RECT 2620.730 1006.090 2621.910 1007.270 ;
        RECT 2619.130 1004.490 2620.310 1005.670 ;
        RECT 2620.730 1004.490 2621.910 1005.670 ;
        RECT 2619.130 826.090 2620.310 827.270 ;
        RECT 2620.730 826.090 2621.910 827.270 ;
        RECT 2619.130 824.490 2620.310 825.670 ;
        RECT 2620.730 824.490 2621.910 825.670 ;
        RECT 2619.130 646.090 2620.310 647.270 ;
        RECT 2620.730 646.090 2621.910 647.270 ;
        RECT 2619.130 644.490 2620.310 645.670 ;
        RECT 2620.730 644.490 2621.910 645.670 ;
        RECT 2619.130 466.090 2620.310 467.270 ;
        RECT 2620.730 466.090 2621.910 467.270 ;
        RECT 2619.130 464.490 2620.310 465.670 ;
        RECT 2620.730 464.490 2621.910 465.670 ;
        RECT 2619.130 286.090 2620.310 287.270 ;
        RECT 2620.730 286.090 2621.910 287.270 ;
        RECT 2619.130 284.490 2620.310 285.670 ;
        RECT 2620.730 284.490 2621.910 285.670 ;
        RECT 2619.130 106.090 2620.310 107.270 ;
        RECT 2620.730 106.090 2621.910 107.270 ;
        RECT 2619.130 104.490 2620.310 105.670 ;
        RECT 2620.730 104.490 2621.910 105.670 ;
        RECT 2619.130 -22.110 2620.310 -20.930 ;
        RECT 2620.730 -22.110 2621.910 -20.930 ;
        RECT 2619.130 -23.710 2620.310 -22.530 ;
        RECT 2620.730 -23.710 2621.910 -22.530 ;
        RECT 2799.130 3542.210 2800.310 3543.390 ;
        RECT 2800.730 3542.210 2801.910 3543.390 ;
        RECT 2799.130 3540.610 2800.310 3541.790 ;
        RECT 2800.730 3540.610 2801.910 3541.790 ;
        RECT 2799.130 3346.090 2800.310 3347.270 ;
        RECT 2800.730 3346.090 2801.910 3347.270 ;
        RECT 2799.130 3344.490 2800.310 3345.670 ;
        RECT 2800.730 3344.490 2801.910 3345.670 ;
        RECT 2799.130 3166.090 2800.310 3167.270 ;
        RECT 2800.730 3166.090 2801.910 3167.270 ;
        RECT 2799.130 3164.490 2800.310 3165.670 ;
        RECT 2800.730 3164.490 2801.910 3165.670 ;
        RECT 2799.130 2986.090 2800.310 2987.270 ;
        RECT 2800.730 2986.090 2801.910 2987.270 ;
        RECT 2799.130 2984.490 2800.310 2985.670 ;
        RECT 2800.730 2984.490 2801.910 2985.670 ;
        RECT 2799.130 2806.090 2800.310 2807.270 ;
        RECT 2800.730 2806.090 2801.910 2807.270 ;
        RECT 2799.130 2804.490 2800.310 2805.670 ;
        RECT 2800.730 2804.490 2801.910 2805.670 ;
        RECT 2799.130 2626.090 2800.310 2627.270 ;
        RECT 2800.730 2626.090 2801.910 2627.270 ;
        RECT 2799.130 2624.490 2800.310 2625.670 ;
        RECT 2800.730 2624.490 2801.910 2625.670 ;
        RECT 2799.130 2446.090 2800.310 2447.270 ;
        RECT 2800.730 2446.090 2801.910 2447.270 ;
        RECT 2799.130 2444.490 2800.310 2445.670 ;
        RECT 2800.730 2444.490 2801.910 2445.670 ;
        RECT 2799.130 2266.090 2800.310 2267.270 ;
        RECT 2800.730 2266.090 2801.910 2267.270 ;
        RECT 2799.130 2264.490 2800.310 2265.670 ;
        RECT 2800.730 2264.490 2801.910 2265.670 ;
        RECT 2799.130 2086.090 2800.310 2087.270 ;
        RECT 2800.730 2086.090 2801.910 2087.270 ;
        RECT 2799.130 2084.490 2800.310 2085.670 ;
        RECT 2800.730 2084.490 2801.910 2085.670 ;
        RECT 2799.130 1906.090 2800.310 1907.270 ;
        RECT 2800.730 1906.090 2801.910 1907.270 ;
        RECT 2799.130 1904.490 2800.310 1905.670 ;
        RECT 2800.730 1904.490 2801.910 1905.670 ;
        RECT 2799.130 1726.090 2800.310 1727.270 ;
        RECT 2800.730 1726.090 2801.910 1727.270 ;
        RECT 2799.130 1724.490 2800.310 1725.670 ;
        RECT 2800.730 1724.490 2801.910 1725.670 ;
        RECT 2799.130 1546.090 2800.310 1547.270 ;
        RECT 2800.730 1546.090 2801.910 1547.270 ;
        RECT 2799.130 1544.490 2800.310 1545.670 ;
        RECT 2800.730 1544.490 2801.910 1545.670 ;
        RECT 2799.130 1366.090 2800.310 1367.270 ;
        RECT 2800.730 1366.090 2801.910 1367.270 ;
        RECT 2799.130 1364.490 2800.310 1365.670 ;
        RECT 2800.730 1364.490 2801.910 1365.670 ;
        RECT 2799.130 1186.090 2800.310 1187.270 ;
        RECT 2800.730 1186.090 2801.910 1187.270 ;
        RECT 2799.130 1184.490 2800.310 1185.670 ;
        RECT 2800.730 1184.490 2801.910 1185.670 ;
        RECT 2799.130 1006.090 2800.310 1007.270 ;
        RECT 2800.730 1006.090 2801.910 1007.270 ;
        RECT 2799.130 1004.490 2800.310 1005.670 ;
        RECT 2800.730 1004.490 2801.910 1005.670 ;
        RECT 2799.130 826.090 2800.310 827.270 ;
        RECT 2800.730 826.090 2801.910 827.270 ;
        RECT 2799.130 824.490 2800.310 825.670 ;
        RECT 2800.730 824.490 2801.910 825.670 ;
        RECT 2799.130 646.090 2800.310 647.270 ;
        RECT 2800.730 646.090 2801.910 647.270 ;
        RECT 2799.130 644.490 2800.310 645.670 ;
        RECT 2800.730 644.490 2801.910 645.670 ;
        RECT 2799.130 466.090 2800.310 467.270 ;
        RECT 2800.730 466.090 2801.910 467.270 ;
        RECT 2799.130 464.490 2800.310 465.670 ;
        RECT 2800.730 464.490 2801.910 465.670 ;
        RECT 2799.130 286.090 2800.310 287.270 ;
        RECT 2800.730 286.090 2801.910 287.270 ;
        RECT 2799.130 284.490 2800.310 285.670 ;
        RECT 2800.730 284.490 2801.910 285.670 ;
        RECT 2799.130 106.090 2800.310 107.270 ;
        RECT 2800.730 106.090 2801.910 107.270 ;
        RECT 2799.130 104.490 2800.310 105.670 ;
        RECT 2800.730 104.490 2801.910 105.670 ;
        RECT 2799.130 -22.110 2800.310 -20.930 ;
        RECT 2800.730 -22.110 2801.910 -20.930 ;
        RECT 2799.130 -23.710 2800.310 -22.530 ;
        RECT 2800.730 -23.710 2801.910 -22.530 ;
        RECT 2945.910 3542.210 2947.090 3543.390 ;
        RECT 2947.510 3542.210 2948.690 3543.390 ;
        RECT 2945.910 3540.610 2947.090 3541.790 ;
        RECT 2947.510 3540.610 2948.690 3541.790 ;
        RECT 2945.910 3346.090 2947.090 3347.270 ;
        RECT 2947.510 3346.090 2948.690 3347.270 ;
        RECT 2945.910 3344.490 2947.090 3345.670 ;
        RECT 2947.510 3344.490 2948.690 3345.670 ;
        RECT 2945.910 3166.090 2947.090 3167.270 ;
        RECT 2947.510 3166.090 2948.690 3167.270 ;
        RECT 2945.910 3164.490 2947.090 3165.670 ;
        RECT 2947.510 3164.490 2948.690 3165.670 ;
        RECT 2945.910 2986.090 2947.090 2987.270 ;
        RECT 2947.510 2986.090 2948.690 2987.270 ;
        RECT 2945.910 2984.490 2947.090 2985.670 ;
        RECT 2947.510 2984.490 2948.690 2985.670 ;
        RECT 2945.910 2806.090 2947.090 2807.270 ;
        RECT 2947.510 2806.090 2948.690 2807.270 ;
        RECT 2945.910 2804.490 2947.090 2805.670 ;
        RECT 2947.510 2804.490 2948.690 2805.670 ;
        RECT 2945.910 2626.090 2947.090 2627.270 ;
        RECT 2947.510 2626.090 2948.690 2627.270 ;
        RECT 2945.910 2624.490 2947.090 2625.670 ;
        RECT 2947.510 2624.490 2948.690 2625.670 ;
        RECT 2945.910 2446.090 2947.090 2447.270 ;
        RECT 2947.510 2446.090 2948.690 2447.270 ;
        RECT 2945.910 2444.490 2947.090 2445.670 ;
        RECT 2947.510 2444.490 2948.690 2445.670 ;
        RECT 2945.910 2266.090 2947.090 2267.270 ;
        RECT 2947.510 2266.090 2948.690 2267.270 ;
        RECT 2945.910 2264.490 2947.090 2265.670 ;
        RECT 2947.510 2264.490 2948.690 2265.670 ;
        RECT 2945.910 2086.090 2947.090 2087.270 ;
        RECT 2947.510 2086.090 2948.690 2087.270 ;
        RECT 2945.910 2084.490 2947.090 2085.670 ;
        RECT 2947.510 2084.490 2948.690 2085.670 ;
        RECT 2945.910 1906.090 2947.090 1907.270 ;
        RECT 2947.510 1906.090 2948.690 1907.270 ;
        RECT 2945.910 1904.490 2947.090 1905.670 ;
        RECT 2947.510 1904.490 2948.690 1905.670 ;
        RECT 2945.910 1726.090 2947.090 1727.270 ;
        RECT 2947.510 1726.090 2948.690 1727.270 ;
        RECT 2945.910 1724.490 2947.090 1725.670 ;
        RECT 2947.510 1724.490 2948.690 1725.670 ;
        RECT 2945.910 1546.090 2947.090 1547.270 ;
        RECT 2947.510 1546.090 2948.690 1547.270 ;
        RECT 2945.910 1544.490 2947.090 1545.670 ;
        RECT 2947.510 1544.490 2948.690 1545.670 ;
        RECT 2945.910 1366.090 2947.090 1367.270 ;
        RECT 2947.510 1366.090 2948.690 1367.270 ;
        RECT 2945.910 1364.490 2947.090 1365.670 ;
        RECT 2947.510 1364.490 2948.690 1365.670 ;
        RECT 2945.910 1186.090 2947.090 1187.270 ;
        RECT 2947.510 1186.090 2948.690 1187.270 ;
        RECT 2945.910 1184.490 2947.090 1185.670 ;
        RECT 2947.510 1184.490 2948.690 1185.670 ;
        RECT 2945.910 1006.090 2947.090 1007.270 ;
        RECT 2947.510 1006.090 2948.690 1007.270 ;
        RECT 2945.910 1004.490 2947.090 1005.670 ;
        RECT 2947.510 1004.490 2948.690 1005.670 ;
        RECT 2945.910 826.090 2947.090 827.270 ;
        RECT 2947.510 826.090 2948.690 827.270 ;
        RECT 2945.910 824.490 2947.090 825.670 ;
        RECT 2947.510 824.490 2948.690 825.670 ;
        RECT 2945.910 646.090 2947.090 647.270 ;
        RECT 2947.510 646.090 2948.690 647.270 ;
        RECT 2945.910 644.490 2947.090 645.670 ;
        RECT 2947.510 644.490 2948.690 645.670 ;
        RECT 2945.910 466.090 2947.090 467.270 ;
        RECT 2947.510 466.090 2948.690 467.270 ;
        RECT 2945.910 464.490 2947.090 465.670 ;
        RECT 2947.510 464.490 2948.690 465.670 ;
        RECT 2945.910 286.090 2947.090 287.270 ;
        RECT 2947.510 286.090 2948.690 287.270 ;
        RECT 2945.910 284.490 2947.090 285.670 ;
        RECT 2947.510 284.490 2948.690 285.670 ;
        RECT 2945.910 106.090 2947.090 107.270 ;
        RECT 2947.510 106.090 2948.690 107.270 ;
        RECT 2945.910 104.490 2947.090 105.670 ;
        RECT 2947.510 104.490 2948.690 105.670 ;
        RECT 2945.910 -22.110 2947.090 -20.930 ;
        RECT 2947.510 -22.110 2948.690 -20.930 ;
        RECT 2945.910 -23.710 2947.090 -22.530 ;
        RECT 2947.510 -23.710 2948.690 -22.530 ;
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
        RECT -43.630 3344.330 2963.250 3347.430 ;
        RECT -43.630 3164.330 2963.250 3167.430 ;
        RECT -43.630 2984.330 2963.250 2987.430 ;
        RECT -43.630 2804.330 2963.250 2807.430 ;
        RECT -43.630 2624.330 2963.250 2627.430 ;
        RECT -43.630 2444.330 2963.250 2447.430 ;
        RECT -43.630 2264.330 2963.250 2267.430 ;
        RECT -43.630 2084.330 2963.250 2087.430 ;
        RECT -43.630 1904.330 2963.250 1907.430 ;
        RECT -43.630 1724.330 2963.250 1727.430 ;
        RECT -43.630 1544.330 2963.250 1547.430 ;
        RECT -43.630 1364.330 2963.250 1367.430 ;
        RECT -43.630 1184.330 2963.250 1187.430 ;
        RECT -43.630 1004.330 2963.250 1007.430 ;
        RECT -43.630 824.330 2963.250 827.430 ;
        RECT -43.630 644.330 2963.250 647.430 ;
        RECT -43.630 464.330 2963.250 467.430 ;
        RECT -43.630 284.330 2963.250 287.430 ;
        RECT -43.630 104.330 2963.250 107.430 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
        RECT 143.970 -38.270 147.070 3557.950 ;
        RECT 323.970 -38.270 327.070 3557.950 ;
        RECT 503.970 810.000 507.070 3557.950 ;
        RECT 683.970 810.000 687.070 3557.950 ;
        RECT 503.970 -38.270 507.070 490.000 ;
        RECT 683.970 -38.270 687.070 490.000 ;
        RECT 863.970 -38.270 867.070 3557.950 ;
        RECT 1043.970 -38.270 1047.070 3557.950 ;
        RECT 1223.970 -38.270 1227.070 3557.950 ;
        RECT 1403.970 -38.270 1407.070 3557.950 ;
        RECT 1583.970 -38.270 1587.070 3557.950 ;
        RECT 1763.970 -38.270 1767.070 3557.950 ;
        RECT 1943.970 -38.270 1947.070 3557.950 ;
        RECT 2123.970 -38.270 2127.070 3557.950 ;
        RECT 2303.970 -38.270 2307.070 3557.950 ;
        RECT 2483.970 -38.270 2487.070 3557.950 ;
        RECT 2663.970 -38.270 2667.070 3557.950 ;
        RECT 2843.970 -38.270 2847.070 3557.950 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
      LAYER via4 ;
        RECT -38.670 3551.810 -37.490 3552.990 ;
        RECT -37.070 3551.810 -35.890 3552.990 ;
        RECT -38.670 3550.210 -37.490 3551.390 ;
        RECT -37.070 3550.210 -35.890 3551.390 ;
        RECT -38.670 3391.090 -37.490 3392.270 ;
        RECT -37.070 3391.090 -35.890 3392.270 ;
        RECT -38.670 3389.490 -37.490 3390.670 ;
        RECT -37.070 3389.490 -35.890 3390.670 ;
        RECT -38.670 3211.090 -37.490 3212.270 ;
        RECT -37.070 3211.090 -35.890 3212.270 ;
        RECT -38.670 3209.490 -37.490 3210.670 ;
        RECT -37.070 3209.490 -35.890 3210.670 ;
        RECT -38.670 3031.090 -37.490 3032.270 ;
        RECT -37.070 3031.090 -35.890 3032.270 ;
        RECT -38.670 3029.490 -37.490 3030.670 ;
        RECT -37.070 3029.490 -35.890 3030.670 ;
        RECT -38.670 2851.090 -37.490 2852.270 ;
        RECT -37.070 2851.090 -35.890 2852.270 ;
        RECT -38.670 2849.490 -37.490 2850.670 ;
        RECT -37.070 2849.490 -35.890 2850.670 ;
        RECT -38.670 2671.090 -37.490 2672.270 ;
        RECT -37.070 2671.090 -35.890 2672.270 ;
        RECT -38.670 2669.490 -37.490 2670.670 ;
        RECT -37.070 2669.490 -35.890 2670.670 ;
        RECT -38.670 2491.090 -37.490 2492.270 ;
        RECT -37.070 2491.090 -35.890 2492.270 ;
        RECT -38.670 2489.490 -37.490 2490.670 ;
        RECT -37.070 2489.490 -35.890 2490.670 ;
        RECT -38.670 2311.090 -37.490 2312.270 ;
        RECT -37.070 2311.090 -35.890 2312.270 ;
        RECT -38.670 2309.490 -37.490 2310.670 ;
        RECT -37.070 2309.490 -35.890 2310.670 ;
        RECT -38.670 2131.090 -37.490 2132.270 ;
        RECT -37.070 2131.090 -35.890 2132.270 ;
        RECT -38.670 2129.490 -37.490 2130.670 ;
        RECT -37.070 2129.490 -35.890 2130.670 ;
        RECT -38.670 1951.090 -37.490 1952.270 ;
        RECT -37.070 1951.090 -35.890 1952.270 ;
        RECT -38.670 1949.490 -37.490 1950.670 ;
        RECT -37.070 1949.490 -35.890 1950.670 ;
        RECT -38.670 1771.090 -37.490 1772.270 ;
        RECT -37.070 1771.090 -35.890 1772.270 ;
        RECT -38.670 1769.490 -37.490 1770.670 ;
        RECT -37.070 1769.490 -35.890 1770.670 ;
        RECT -38.670 1591.090 -37.490 1592.270 ;
        RECT -37.070 1591.090 -35.890 1592.270 ;
        RECT -38.670 1589.490 -37.490 1590.670 ;
        RECT -37.070 1589.490 -35.890 1590.670 ;
        RECT -38.670 1411.090 -37.490 1412.270 ;
        RECT -37.070 1411.090 -35.890 1412.270 ;
        RECT -38.670 1409.490 -37.490 1410.670 ;
        RECT -37.070 1409.490 -35.890 1410.670 ;
        RECT -38.670 1231.090 -37.490 1232.270 ;
        RECT -37.070 1231.090 -35.890 1232.270 ;
        RECT -38.670 1229.490 -37.490 1230.670 ;
        RECT -37.070 1229.490 -35.890 1230.670 ;
        RECT -38.670 1051.090 -37.490 1052.270 ;
        RECT -37.070 1051.090 -35.890 1052.270 ;
        RECT -38.670 1049.490 -37.490 1050.670 ;
        RECT -37.070 1049.490 -35.890 1050.670 ;
        RECT -38.670 871.090 -37.490 872.270 ;
        RECT -37.070 871.090 -35.890 872.270 ;
        RECT -38.670 869.490 -37.490 870.670 ;
        RECT -37.070 869.490 -35.890 870.670 ;
        RECT -38.670 691.090 -37.490 692.270 ;
        RECT -37.070 691.090 -35.890 692.270 ;
        RECT -38.670 689.490 -37.490 690.670 ;
        RECT -37.070 689.490 -35.890 690.670 ;
        RECT -38.670 511.090 -37.490 512.270 ;
        RECT -37.070 511.090 -35.890 512.270 ;
        RECT -38.670 509.490 -37.490 510.670 ;
        RECT -37.070 509.490 -35.890 510.670 ;
        RECT -38.670 331.090 -37.490 332.270 ;
        RECT -37.070 331.090 -35.890 332.270 ;
        RECT -38.670 329.490 -37.490 330.670 ;
        RECT -37.070 329.490 -35.890 330.670 ;
        RECT -38.670 151.090 -37.490 152.270 ;
        RECT -37.070 151.090 -35.890 152.270 ;
        RECT -38.670 149.490 -37.490 150.670 ;
        RECT -37.070 149.490 -35.890 150.670 ;
        RECT -38.670 -31.710 -37.490 -30.530 ;
        RECT -37.070 -31.710 -35.890 -30.530 ;
        RECT -38.670 -33.310 -37.490 -32.130 ;
        RECT -37.070 -33.310 -35.890 -32.130 ;
        RECT 144.130 3551.810 145.310 3552.990 ;
        RECT 145.730 3551.810 146.910 3552.990 ;
        RECT 144.130 3550.210 145.310 3551.390 ;
        RECT 145.730 3550.210 146.910 3551.390 ;
        RECT 144.130 3391.090 145.310 3392.270 ;
        RECT 145.730 3391.090 146.910 3392.270 ;
        RECT 144.130 3389.490 145.310 3390.670 ;
        RECT 145.730 3389.490 146.910 3390.670 ;
        RECT 144.130 3211.090 145.310 3212.270 ;
        RECT 145.730 3211.090 146.910 3212.270 ;
        RECT 144.130 3209.490 145.310 3210.670 ;
        RECT 145.730 3209.490 146.910 3210.670 ;
        RECT 144.130 3031.090 145.310 3032.270 ;
        RECT 145.730 3031.090 146.910 3032.270 ;
        RECT 144.130 3029.490 145.310 3030.670 ;
        RECT 145.730 3029.490 146.910 3030.670 ;
        RECT 144.130 2851.090 145.310 2852.270 ;
        RECT 145.730 2851.090 146.910 2852.270 ;
        RECT 144.130 2849.490 145.310 2850.670 ;
        RECT 145.730 2849.490 146.910 2850.670 ;
        RECT 144.130 2671.090 145.310 2672.270 ;
        RECT 145.730 2671.090 146.910 2672.270 ;
        RECT 144.130 2669.490 145.310 2670.670 ;
        RECT 145.730 2669.490 146.910 2670.670 ;
        RECT 144.130 2491.090 145.310 2492.270 ;
        RECT 145.730 2491.090 146.910 2492.270 ;
        RECT 144.130 2489.490 145.310 2490.670 ;
        RECT 145.730 2489.490 146.910 2490.670 ;
        RECT 144.130 2311.090 145.310 2312.270 ;
        RECT 145.730 2311.090 146.910 2312.270 ;
        RECT 144.130 2309.490 145.310 2310.670 ;
        RECT 145.730 2309.490 146.910 2310.670 ;
        RECT 144.130 2131.090 145.310 2132.270 ;
        RECT 145.730 2131.090 146.910 2132.270 ;
        RECT 144.130 2129.490 145.310 2130.670 ;
        RECT 145.730 2129.490 146.910 2130.670 ;
        RECT 144.130 1951.090 145.310 1952.270 ;
        RECT 145.730 1951.090 146.910 1952.270 ;
        RECT 144.130 1949.490 145.310 1950.670 ;
        RECT 145.730 1949.490 146.910 1950.670 ;
        RECT 144.130 1771.090 145.310 1772.270 ;
        RECT 145.730 1771.090 146.910 1772.270 ;
        RECT 144.130 1769.490 145.310 1770.670 ;
        RECT 145.730 1769.490 146.910 1770.670 ;
        RECT 144.130 1591.090 145.310 1592.270 ;
        RECT 145.730 1591.090 146.910 1592.270 ;
        RECT 144.130 1589.490 145.310 1590.670 ;
        RECT 145.730 1589.490 146.910 1590.670 ;
        RECT 144.130 1411.090 145.310 1412.270 ;
        RECT 145.730 1411.090 146.910 1412.270 ;
        RECT 144.130 1409.490 145.310 1410.670 ;
        RECT 145.730 1409.490 146.910 1410.670 ;
        RECT 144.130 1231.090 145.310 1232.270 ;
        RECT 145.730 1231.090 146.910 1232.270 ;
        RECT 144.130 1229.490 145.310 1230.670 ;
        RECT 145.730 1229.490 146.910 1230.670 ;
        RECT 144.130 1051.090 145.310 1052.270 ;
        RECT 145.730 1051.090 146.910 1052.270 ;
        RECT 144.130 1049.490 145.310 1050.670 ;
        RECT 145.730 1049.490 146.910 1050.670 ;
        RECT 144.130 871.090 145.310 872.270 ;
        RECT 145.730 871.090 146.910 872.270 ;
        RECT 144.130 869.490 145.310 870.670 ;
        RECT 145.730 869.490 146.910 870.670 ;
        RECT 144.130 691.090 145.310 692.270 ;
        RECT 145.730 691.090 146.910 692.270 ;
        RECT 144.130 689.490 145.310 690.670 ;
        RECT 145.730 689.490 146.910 690.670 ;
        RECT 144.130 511.090 145.310 512.270 ;
        RECT 145.730 511.090 146.910 512.270 ;
        RECT 144.130 509.490 145.310 510.670 ;
        RECT 145.730 509.490 146.910 510.670 ;
        RECT 144.130 331.090 145.310 332.270 ;
        RECT 145.730 331.090 146.910 332.270 ;
        RECT 144.130 329.490 145.310 330.670 ;
        RECT 145.730 329.490 146.910 330.670 ;
        RECT 144.130 151.090 145.310 152.270 ;
        RECT 145.730 151.090 146.910 152.270 ;
        RECT 144.130 149.490 145.310 150.670 ;
        RECT 145.730 149.490 146.910 150.670 ;
        RECT 144.130 -31.710 145.310 -30.530 ;
        RECT 145.730 -31.710 146.910 -30.530 ;
        RECT 144.130 -33.310 145.310 -32.130 ;
        RECT 145.730 -33.310 146.910 -32.130 ;
        RECT 324.130 3551.810 325.310 3552.990 ;
        RECT 325.730 3551.810 326.910 3552.990 ;
        RECT 324.130 3550.210 325.310 3551.390 ;
        RECT 325.730 3550.210 326.910 3551.390 ;
        RECT 324.130 3391.090 325.310 3392.270 ;
        RECT 325.730 3391.090 326.910 3392.270 ;
        RECT 324.130 3389.490 325.310 3390.670 ;
        RECT 325.730 3389.490 326.910 3390.670 ;
        RECT 324.130 3211.090 325.310 3212.270 ;
        RECT 325.730 3211.090 326.910 3212.270 ;
        RECT 324.130 3209.490 325.310 3210.670 ;
        RECT 325.730 3209.490 326.910 3210.670 ;
        RECT 324.130 3031.090 325.310 3032.270 ;
        RECT 325.730 3031.090 326.910 3032.270 ;
        RECT 324.130 3029.490 325.310 3030.670 ;
        RECT 325.730 3029.490 326.910 3030.670 ;
        RECT 324.130 2851.090 325.310 2852.270 ;
        RECT 325.730 2851.090 326.910 2852.270 ;
        RECT 324.130 2849.490 325.310 2850.670 ;
        RECT 325.730 2849.490 326.910 2850.670 ;
        RECT 324.130 2671.090 325.310 2672.270 ;
        RECT 325.730 2671.090 326.910 2672.270 ;
        RECT 324.130 2669.490 325.310 2670.670 ;
        RECT 325.730 2669.490 326.910 2670.670 ;
        RECT 324.130 2491.090 325.310 2492.270 ;
        RECT 325.730 2491.090 326.910 2492.270 ;
        RECT 324.130 2489.490 325.310 2490.670 ;
        RECT 325.730 2489.490 326.910 2490.670 ;
        RECT 324.130 2311.090 325.310 2312.270 ;
        RECT 325.730 2311.090 326.910 2312.270 ;
        RECT 324.130 2309.490 325.310 2310.670 ;
        RECT 325.730 2309.490 326.910 2310.670 ;
        RECT 324.130 2131.090 325.310 2132.270 ;
        RECT 325.730 2131.090 326.910 2132.270 ;
        RECT 324.130 2129.490 325.310 2130.670 ;
        RECT 325.730 2129.490 326.910 2130.670 ;
        RECT 324.130 1951.090 325.310 1952.270 ;
        RECT 325.730 1951.090 326.910 1952.270 ;
        RECT 324.130 1949.490 325.310 1950.670 ;
        RECT 325.730 1949.490 326.910 1950.670 ;
        RECT 324.130 1771.090 325.310 1772.270 ;
        RECT 325.730 1771.090 326.910 1772.270 ;
        RECT 324.130 1769.490 325.310 1770.670 ;
        RECT 325.730 1769.490 326.910 1770.670 ;
        RECT 324.130 1591.090 325.310 1592.270 ;
        RECT 325.730 1591.090 326.910 1592.270 ;
        RECT 324.130 1589.490 325.310 1590.670 ;
        RECT 325.730 1589.490 326.910 1590.670 ;
        RECT 324.130 1411.090 325.310 1412.270 ;
        RECT 325.730 1411.090 326.910 1412.270 ;
        RECT 324.130 1409.490 325.310 1410.670 ;
        RECT 325.730 1409.490 326.910 1410.670 ;
        RECT 324.130 1231.090 325.310 1232.270 ;
        RECT 325.730 1231.090 326.910 1232.270 ;
        RECT 324.130 1229.490 325.310 1230.670 ;
        RECT 325.730 1229.490 326.910 1230.670 ;
        RECT 324.130 1051.090 325.310 1052.270 ;
        RECT 325.730 1051.090 326.910 1052.270 ;
        RECT 324.130 1049.490 325.310 1050.670 ;
        RECT 325.730 1049.490 326.910 1050.670 ;
        RECT 324.130 871.090 325.310 872.270 ;
        RECT 325.730 871.090 326.910 872.270 ;
        RECT 324.130 869.490 325.310 870.670 ;
        RECT 325.730 869.490 326.910 870.670 ;
        RECT 504.130 3551.810 505.310 3552.990 ;
        RECT 505.730 3551.810 506.910 3552.990 ;
        RECT 504.130 3550.210 505.310 3551.390 ;
        RECT 505.730 3550.210 506.910 3551.390 ;
        RECT 504.130 3391.090 505.310 3392.270 ;
        RECT 505.730 3391.090 506.910 3392.270 ;
        RECT 504.130 3389.490 505.310 3390.670 ;
        RECT 505.730 3389.490 506.910 3390.670 ;
        RECT 504.130 3211.090 505.310 3212.270 ;
        RECT 505.730 3211.090 506.910 3212.270 ;
        RECT 504.130 3209.490 505.310 3210.670 ;
        RECT 505.730 3209.490 506.910 3210.670 ;
        RECT 504.130 3031.090 505.310 3032.270 ;
        RECT 505.730 3031.090 506.910 3032.270 ;
        RECT 504.130 3029.490 505.310 3030.670 ;
        RECT 505.730 3029.490 506.910 3030.670 ;
        RECT 504.130 2851.090 505.310 2852.270 ;
        RECT 505.730 2851.090 506.910 2852.270 ;
        RECT 504.130 2849.490 505.310 2850.670 ;
        RECT 505.730 2849.490 506.910 2850.670 ;
        RECT 504.130 2671.090 505.310 2672.270 ;
        RECT 505.730 2671.090 506.910 2672.270 ;
        RECT 504.130 2669.490 505.310 2670.670 ;
        RECT 505.730 2669.490 506.910 2670.670 ;
        RECT 504.130 2491.090 505.310 2492.270 ;
        RECT 505.730 2491.090 506.910 2492.270 ;
        RECT 504.130 2489.490 505.310 2490.670 ;
        RECT 505.730 2489.490 506.910 2490.670 ;
        RECT 504.130 2311.090 505.310 2312.270 ;
        RECT 505.730 2311.090 506.910 2312.270 ;
        RECT 504.130 2309.490 505.310 2310.670 ;
        RECT 505.730 2309.490 506.910 2310.670 ;
        RECT 504.130 2131.090 505.310 2132.270 ;
        RECT 505.730 2131.090 506.910 2132.270 ;
        RECT 504.130 2129.490 505.310 2130.670 ;
        RECT 505.730 2129.490 506.910 2130.670 ;
        RECT 504.130 1951.090 505.310 1952.270 ;
        RECT 505.730 1951.090 506.910 1952.270 ;
        RECT 504.130 1949.490 505.310 1950.670 ;
        RECT 505.730 1949.490 506.910 1950.670 ;
        RECT 504.130 1771.090 505.310 1772.270 ;
        RECT 505.730 1771.090 506.910 1772.270 ;
        RECT 504.130 1769.490 505.310 1770.670 ;
        RECT 505.730 1769.490 506.910 1770.670 ;
        RECT 504.130 1591.090 505.310 1592.270 ;
        RECT 505.730 1591.090 506.910 1592.270 ;
        RECT 504.130 1589.490 505.310 1590.670 ;
        RECT 505.730 1589.490 506.910 1590.670 ;
        RECT 504.130 1411.090 505.310 1412.270 ;
        RECT 505.730 1411.090 506.910 1412.270 ;
        RECT 504.130 1409.490 505.310 1410.670 ;
        RECT 505.730 1409.490 506.910 1410.670 ;
        RECT 504.130 1231.090 505.310 1232.270 ;
        RECT 505.730 1231.090 506.910 1232.270 ;
        RECT 504.130 1229.490 505.310 1230.670 ;
        RECT 505.730 1229.490 506.910 1230.670 ;
        RECT 504.130 1051.090 505.310 1052.270 ;
        RECT 505.730 1051.090 506.910 1052.270 ;
        RECT 504.130 1049.490 505.310 1050.670 ;
        RECT 505.730 1049.490 506.910 1050.670 ;
        RECT 504.130 871.090 505.310 872.270 ;
        RECT 505.730 871.090 506.910 872.270 ;
        RECT 504.130 869.490 505.310 870.670 ;
        RECT 505.730 869.490 506.910 870.670 ;
        RECT 684.130 3551.810 685.310 3552.990 ;
        RECT 685.730 3551.810 686.910 3552.990 ;
        RECT 684.130 3550.210 685.310 3551.390 ;
        RECT 685.730 3550.210 686.910 3551.390 ;
        RECT 684.130 3391.090 685.310 3392.270 ;
        RECT 685.730 3391.090 686.910 3392.270 ;
        RECT 684.130 3389.490 685.310 3390.670 ;
        RECT 685.730 3389.490 686.910 3390.670 ;
        RECT 684.130 3211.090 685.310 3212.270 ;
        RECT 685.730 3211.090 686.910 3212.270 ;
        RECT 684.130 3209.490 685.310 3210.670 ;
        RECT 685.730 3209.490 686.910 3210.670 ;
        RECT 684.130 3031.090 685.310 3032.270 ;
        RECT 685.730 3031.090 686.910 3032.270 ;
        RECT 684.130 3029.490 685.310 3030.670 ;
        RECT 685.730 3029.490 686.910 3030.670 ;
        RECT 684.130 2851.090 685.310 2852.270 ;
        RECT 685.730 2851.090 686.910 2852.270 ;
        RECT 684.130 2849.490 685.310 2850.670 ;
        RECT 685.730 2849.490 686.910 2850.670 ;
        RECT 684.130 2671.090 685.310 2672.270 ;
        RECT 685.730 2671.090 686.910 2672.270 ;
        RECT 684.130 2669.490 685.310 2670.670 ;
        RECT 685.730 2669.490 686.910 2670.670 ;
        RECT 684.130 2491.090 685.310 2492.270 ;
        RECT 685.730 2491.090 686.910 2492.270 ;
        RECT 684.130 2489.490 685.310 2490.670 ;
        RECT 685.730 2489.490 686.910 2490.670 ;
        RECT 684.130 2311.090 685.310 2312.270 ;
        RECT 685.730 2311.090 686.910 2312.270 ;
        RECT 684.130 2309.490 685.310 2310.670 ;
        RECT 685.730 2309.490 686.910 2310.670 ;
        RECT 684.130 2131.090 685.310 2132.270 ;
        RECT 685.730 2131.090 686.910 2132.270 ;
        RECT 684.130 2129.490 685.310 2130.670 ;
        RECT 685.730 2129.490 686.910 2130.670 ;
        RECT 684.130 1951.090 685.310 1952.270 ;
        RECT 685.730 1951.090 686.910 1952.270 ;
        RECT 684.130 1949.490 685.310 1950.670 ;
        RECT 685.730 1949.490 686.910 1950.670 ;
        RECT 684.130 1771.090 685.310 1772.270 ;
        RECT 685.730 1771.090 686.910 1772.270 ;
        RECT 684.130 1769.490 685.310 1770.670 ;
        RECT 685.730 1769.490 686.910 1770.670 ;
        RECT 684.130 1591.090 685.310 1592.270 ;
        RECT 685.730 1591.090 686.910 1592.270 ;
        RECT 684.130 1589.490 685.310 1590.670 ;
        RECT 685.730 1589.490 686.910 1590.670 ;
        RECT 684.130 1411.090 685.310 1412.270 ;
        RECT 685.730 1411.090 686.910 1412.270 ;
        RECT 684.130 1409.490 685.310 1410.670 ;
        RECT 685.730 1409.490 686.910 1410.670 ;
        RECT 684.130 1231.090 685.310 1232.270 ;
        RECT 685.730 1231.090 686.910 1232.270 ;
        RECT 684.130 1229.490 685.310 1230.670 ;
        RECT 685.730 1229.490 686.910 1230.670 ;
        RECT 684.130 1051.090 685.310 1052.270 ;
        RECT 685.730 1051.090 686.910 1052.270 ;
        RECT 684.130 1049.490 685.310 1050.670 ;
        RECT 685.730 1049.490 686.910 1050.670 ;
        RECT 684.130 871.090 685.310 872.270 ;
        RECT 685.730 871.090 686.910 872.270 ;
        RECT 684.130 869.490 685.310 870.670 ;
        RECT 685.730 869.490 686.910 870.670 ;
        RECT 864.130 3551.810 865.310 3552.990 ;
        RECT 865.730 3551.810 866.910 3552.990 ;
        RECT 864.130 3550.210 865.310 3551.390 ;
        RECT 865.730 3550.210 866.910 3551.390 ;
        RECT 864.130 3391.090 865.310 3392.270 ;
        RECT 865.730 3391.090 866.910 3392.270 ;
        RECT 864.130 3389.490 865.310 3390.670 ;
        RECT 865.730 3389.490 866.910 3390.670 ;
        RECT 864.130 3211.090 865.310 3212.270 ;
        RECT 865.730 3211.090 866.910 3212.270 ;
        RECT 864.130 3209.490 865.310 3210.670 ;
        RECT 865.730 3209.490 866.910 3210.670 ;
        RECT 864.130 3031.090 865.310 3032.270 ;
        RECT 865.730 3031.090 866.910 3032.270 ;
        RECT 864.130 3029.490 865.310 3030.670 ;
        RECT 865.730 3029.490 866.910 3030.670 ;
        RECT 864.130 2851.090 865.310 2852.270 ;
        RECT 865.730 2851.090 866.910 2852.270 ;
        RECT 864.130 2849.490 865.310 2850.670 ;
        RECT 865.730 2849.490 866.910 2850.670 ;
        RECT 864.130 2671.090 865.310 2672.270 ;
        RECT 865.730 2671.090 866.910 2672.270 ;
        RECT 864.130 2669.490 865.310 2670.670 ;
        RECT 865.730 2669.490 866.910 2670.670 ;
        RECT 864.130 2491.090 865.310 2492.270 ;
        RECT 865.730 2491.090 866.910 2492.270 ;
        RECT 864.130 2489.490 865.310 2490.670 ;
        RECT 865.730 2489.490 866.910 2490.670 ;
        RECT 864.130 2311.090 865.310 2312.270 ;
        RECT 865.730 2311.090 866.910 2312.270 ;
        RECT 864.130 2309.490 865.310 2310.670 ;
        RECT 865.730 2309.490 866.910 2310.670 ;
        RECT 864.130 2131.090 865.310 2132.270 ;
        RECT 865.730 2131.090 866.910 2132.270 ;
        RECT 864.130 2129.490 865.310 2130.670 ;
        RECT 865.730 2129.490 866.910 2130.670 ;
        RECT 864.130 1951.090 865.310 1952.270 ;
        RECT 865.730 1951.090 866.910 1952.270 ;
        RECT 864.130 1949.490 865.310 1950.670 ;
        RECT 865.730 1949.490 866.910 1950.670 ;
        RECT 864.130 1771.090 865.310 1772.270 ;
        RECT 865.730 1771.090 866.910 1772.270 ;
        RECT 864.130 1769.490 865.310 1770.670 ;
        RECT 865.730 1769.490 866.910 1770.670 ;
        RECT 864.130 1591.090 865.310 1592.270 ;
        RECT 865.730 1591.090 866.910 1592.270 ;
        RECT 864.130 1589.490 865.310 1590.670 ;
        RECT 865.730 1589.490 866.910 1590.670 ;
        RECT 864.130 1411.090 865.310 1412.270 ;
        RECT 865.730 1411.090 866.910 1412.270 ;
        RECT 864.130 1409.490 865.310 1410.670 ;
        RECT 865.730 1409.490 866.910 1410.670 ;
        RECT 864.130 1231.090 865.310 1232.270 ;
        RECT 865.730 1231.090 866.910 1232.270 ;
        RECT 864.130 1229.490 865.310 1230.670 ;
        RECT 865.730 1229.490 866.910 1230.670 ;
        RECT 864.130 1051.090 865.310 1052.270 ;
        RECT 865.730 1051.090 866.910 1052.270 ;
        RECT 864.130 1049.490 865.310 1050.670 ;
        RECT 865.730 1049.490 866.910 1050.670 ;
        RECT 864.130 871.090 865.310 872.270 ;
        RECT 865.730 871.090 866.910 872.270 ;
        RECT 864.130 869.490 865.310 870.670 ;
        RECT 865.730 869.490 866.910 870.670 ;
        RECT 324.130 691.090 325.310 692.270 ;
        RECT 325.730 691.090 326.910 692.270 ;
        RECT 324.130 689.490 325.310 690.670 ;
        RECT 325.730 689.490 326.910 690.670 ;
        RECT 324.130 511.090 325.310 512.270 ;
        RECT 325.730 511.090 326.910 512.270 ;
        RECT 324.130 509.490 325.310 510.670 ;
        RECT 325.730 509.490 326.910 510.670 ;
        RECT 864.130 691.090 865.310 692.270 ;
        RECT 865.730 691.090 866.910 692.270 ;
        RECT 864.130 689.490 865.310 690.670 ;
        RECT 865.730 689.490 866.910 690.670 ;
        RECT 864.130 511.090 865.310 512.270 ;
        RECT 865.730 511.090 866.910 512.270 ;
        RECT 864.130 509.490 865.310 510.670 ;
        RECT 865.730 509.490 866.910 510.670 ;
        RECT 324.130 331.090 325.310 332.270 ;
        RECT 325.730 331.090 326.910 332.270 ;
        RECT 324.130 329.490 325.310 330.670 ;
        RECT 325.730 329.490 326.910 330.670 ;
        RECT 324.130 151.090 325.310 152.270 ;
        RECT 325.730 151.090 326.910 152.270 ;
        RECT 324.130 149.490 325.310 150.670 ;
        RECT 325.730 149.490 326.910 150.670 ;
        RECT 324.130 -31.710 325.310 -30.530 ;
        RECT 325.730 -31.710 326.910 -30.530 ;
        RECT 324.130 -33.310 325.310 -32.130 ;
        RECT 325.730 -33.310 326.910 -32.130 ;
        RECT 504.130 331.090 505.310 332.270 ;
        RECT 505.730 331.090 506.910 332.270 ;
        RECT 504.130 329.490 505.310 330.670 ;
        RECT 505.730 329.490 506.910 330.670 ;
        RECT 504.130 151.090 505.310 152.270 ;
        RECT 505.730 151.090 506.910 152.270 ;
        RECT 504.130 149.490 505.310 150.670 ;
        RECT 505.730 149.490 506.910 150.670 ;
        RECT 504.130 -31.710 505.310 -30.530 ;
        RECT 505.730 -31.710 506.910 -30.530 ;
        RECT 504.130 -33.310 505.310 -32.130 ;
        RECT 505.730 -33.310 506.910 -32.130 ;
        RECT 684.130 331.090 685.310 332.270 ;
        RECT 685.730 331.090 686.910 332.270 ;
        RECT 684.130 329.490 685.310 330.670 ;
        RECT 685.730 329.490 686.910 330.670 ;
        RECT 684.130 151.090 685.310 152.270 ;
        RECT 685.730 151.090 686.910 152.270 ;
        RECT 684.130 149.490 685.310 150.670 ;
        RECT 685.730 149.490 686.910 150.670 ;
        RECT 684.130 -31.710 685.310 -30.530 ;
        RECT 685.730 -31.710 686.910 -30.530 ;
        RECT 684.130 -33.310 685.310 -32.130 ;
        RECT 685.730 -33.310 686.910 -32.130 ;
        RECT 864.130 331.090 865.310 332.270 ;
        RECT 865.730 331.090 866.910 332.270 ;
        RECT 864.130 329.490 865.310 330.670 ;
        RECT 865.730 329.490 866.910 330.670 ;
        RECT 864.130 151.090 865.310 152.270 ;
        RECT 865.730 151.090 866.910 152.270 ;
        RECT 864.130 149.490 865.310 150.670 ;
        RECT 865.730 149.490 866.910 150.670 ;
        RECT 864.130 -31.710 865.310 -30.530 ;
        RECT 865.730 -31.710 866.910 -30.530 ;
        RECT 864.130 -33.310 865.310 -32.130 ;
        RECT 865.730 -33.310 866.910 -32.130 ;
        RECT 1044.130 3551.810 1045.310 3552.990 ;
        RECT 1045.730 3551.810 1046.910 3552.990 ;
        RECT 1044.130 3550.210 1045.310 3551.390 ;
        RECT 1045.730 3550.210 1046.910 3551.390 ;
        RECT 1044.130 3391.090 1045.310 3392.270 ;
        RECT 1045.730 3391.090 1046.910 3392.270 ;
        RECT 1044.130 3389.490 1045.310 3390.670 ;
        RECT 1045.730 3389.490 1046.910 3390.670 ;
        RECT 1044.130 3211.090 1045.310 3212.270 ;
        RECT 1045.730 3211.090 1046.910 3212.270 ;
        RECT 1044.130 3209.490 1045.310 3210.670 ;
        RECT 1045.730 3209.490 1046.910 3210.670 ;
        RECT 1044.130 3031.090 1045.310 3032.270 ;
        RECT 1045.730 3031.090 1046.910 3032.270 ;
        RECT 1044.130 3029.490 1045.310 3030.670 ;
        RECT 1045.730 3029.490 1046.910 3030.670 ;
        RECT 1044.130 2851.090 1045.310 2852.270 ;
        RECT 1045.730 2851.090 1046.910 2852.270 ;
        RECT 1044.130 2849.490 1045.310 2850.670 ;
        RECT 1045.730 2849.490 1046.910 2850.670 ;
        RECT 1044.130 2671.090 1045.310 2672.270 ;
        RECT 1045.730 2671.090 1046.910 2672.270 ;
        RECT 1044.130 2669.490 1045.310 2670.670 ;
        RECT 1045.730 2669.490 1046.910 2670.670 ;
        RECT 1044.130 2491.090 1045.310 2492.270 ;
        RECT 1045.730 2491.090 1046.910 2492.270 ;
        RECT 1044.130 2489.490 1045.310 2490.670 ;
        RECT 1045.730 2489.490 1046.910 2490.670 ;
        RECT 1044.130 2311.090 1045.310 2312.270 ;
        RECT 1045.730 2311.090 1046.910 2312.270 ;
        RECT 1044.130 2309.490 1045.310 2310.670 ;
        RECT 1045.730 2309.490 1046.910 2310.670 ;
        RECT 1044.130 2131.090 1045.310 2132.270 ;
        RECT 1045.730 2131.090 1046.910 2132.270 ;
        RECT 1044.130 2129.490 1045.310 2130.670 ;
        RECT 1045.730 2129.490 1046.910 2130.670 ;
        RECT 1044.130 1951.090 1045.310 1952.270 ;
        RECT 1045.730 1951.090 1046.910 1952.270 ;
        RECT 1044.130 1949.490 1045.310 1950.670 ;
        RECT 1045.730 1949.490 1046.910 1950.670 ;
        RECT 1044.130 1771.090 1045.310 1772.270 ;
        RECT 1045.730 1771.090 1046.910 1772.270 ;
        RECT 1044.130 1769.490 1045.310 1770.670 ;
        RECT 1045.730 1769.490 1046.910 1770.670 ;
        RECT 1044.130 1591.090 1045.310 1592.270 ;
        RECT 1045.730 1591.090 1046.910 1592.270 ;
        RECT 1044.130 1589.490 1045.310 1590.670 ;
        RECT 1045.730 1589.490 1046.910 1590.670 ;
        RECT 1044.130 1411.090 1045.310 1412.270 ;
        RECT 1045.730 1411.090 1046.910 1412.270 ;
        RECT 1044.130 1409.490 1045.310 1410.670 ;
        RECT 1045.730 1409.490 1046.910 1410.670 ;
        RECT 1044.130 1231.090 1045.310 1232.270 ;
        RECT 1045.730 1231.090 1046.910 1232.270 ;
        RECT 1044.130 1229.490 1045.310 1230.670 ;
        RECT 1045.730 1229.490 1046.910 1230.670 ;
        RECT 1044.130 1051.090 1045.310 1052.270 ;
        RECT 1045.730 1051.090 1046.910 1052.270 ;
        RECT 1044.130 1049.490 1045.310 1050.670 ;
        RECT 1045.730 1049.490 1046.910 1050.670 ;
        RECT 1044.130 871.090 1045.310 872.270 ;
        RECT 1045.730 871.090 1046.910 872.270 ;
        RECT 1044.130 869.490 1045.310 870.670 ;
        RECT 1045.730 869.490 1046.910 870.670 ;
        RECT 1044.130 691.090 1045.310 692.270 ;
        RECT 1045.730 691.090 1046.910 692.270 ;
        RECT 1044.130 689.490 1045.310 690.670 ;
        RECT 1045.730 689.490 1046.910 690.670 ;
        RECT 1044.130 511.090 1045.310 512.270 ;
        RECT 1045.730 511.090 1046.910 512.270 ;
        RECT 1044.130 509.490 1045.310 510.670 ;
        RECT 1045.730 509.490 1046.910 510.670 ;
        RECT 1044.130 331.090 1045.310 332.270 ;
        RECT 1045.730 331.090 1046.910 332.270 ;
        RECT 1044.130 329.490 1045.310 330.670 ;
        RECT 1045.730 329.490 1046.910 330.670 ;
        RECT 1044.130 151.090 1045.310 152.270 ;
        RECT 1045.730 151.090 1046.910 152.270 ;
        RECT 1044.130 149.490 1045.310 150.670 ;
        RECT 1045.730 149.490 1046.910 150.670 ;
        RECT 1044.130 -31.710 1045.310 -30.530 ;
        RECT 1045.730 -31.710 1046.910 -30.530 ;
        RECT 1044.130 -33.310 1045.310 -32.130 ;
        RECT 1045.730 -33.310 1046.910 -32.130 ;
        RECT 1224.130 3551.810 1225.310 3552.990 ;
        RECT 1225.730 3551.810 1226.910 3552.990 ;
        RECT 1224.130 3550.210 1225.310 3551.390 ;
        RECT 1225.730 3550.210 1226.910 3551.390 ;
        RECT 1224.130 3391.090 1225.310 3392.270 ;
        RECT 1225.730 3391.090 1226.910 3392.270 ;
        RECT 1224.130 3389.490 1225.310 3390.670 ;
        RECT 1225.730 3389.490 1226.910 3390.670 ;
        RECT 1224.130 3211.090 1225.310 3212.270 ;
        RECT 1225.730 3211.090 1226.910 3212.270 ;
        RECT 1224.130 3209.490 1225.310 3210.670 ;
        RECT 1225.730 3209.490 1226.910 3210.670 ;
        RECT 1224.130 3031.090 1225.310 3032.270 ;
        RECT 1225.730 3031.090 1226.910 3032.270 ;
        RECT 1224.130 3029.490 1225.310 3030.670 ;
        RECT 1225.730 3029.490 1226.910 3030.670 ;
        RECT 1224.130 2851.090 1225.310 2852.270 ;
        RECT 1225.730 2851.090 1226.910 2852.270 ;
        RECT 1224.130 2849.490 1225.310 2850.670 ;
        RECT 1225.730 2849.490 1226.910 2850.670 ;
        RECT 1224.130 2671.090 1225.310 2672.270 ;
        RECT 1225.730 2671.090 1226.910 2672.270 ;
        RECT 1224.130 2669.490 1225.310 2670.670 ;
        RECT 1225.730 2669.490 1226.910 2670.670 ;
        RECT 1224.130 2491.090 1225.310 2492.270 ;
        RECT 1225.730 2491.090 1226.910 2492.270 ;
        RECT 1224.130 2489.490 1225.310 2490.670 ;
        RECT 1225.730 2489.490 1226.910 2490.670 ;
        RECT 1224.130 2311.090 1225.310 2312.270 ;
        RECT 1225.730 2311.090 1226.910 2312.270 ;
        RECT 1224.130 2309.490 1225.310 2310.670 ;
        RECT 1225.730 2309.490 1226.910 2310.670 ;
        RECT 1224.130 2131.090 1225.310 2132.270 ;
        RECT 1225.730 2131.090 1226.910 2132.270 ;
        RECT 1224.130 2129.490 1225.310 2130.670 ;
        RECT 1225.730 2129.490 1226.910 2130.670 ;
        RECT 1224.130 1951.090 1225.310 1952.270 ;
        RECT 1225.730 1951.090 1226.910 1952.270 ;
        RECT 1224.130 1949.490 1225.310 1950.670 ;
        RECT 1225.730 1949.490 1226.910 1950.670 ;
        RECT 1224.130 1771.090 1225.310 1772.270 ;
        RECT 1225.730 1771.090 1226.910 1772.270 ;
        RECT 1224.130 1769.490 1225.310 1770.670 ;
        RECT 1225.730 1769.490 1226.910 1770.670 ;
        RECT 1224.130 1591.090 1225.310 1592.270 ;
        RECT 1225.730 1591.090 1226.910 1592.270 ;
        RECT 1224.130 1589.490 1225.310 1590.670 ;
        RECT 1225.730 1589.490 1226.910 1590.670 ;
        RECT 1224.130 1411.090 1225.310 1412.270 ;
        RECT 1225.730 1411.090 1226.910 1412.270 ;
        RECT 1224.130 1409.490 1225.310 1410.670 ;
        RECT 1225.730 1409.490 1226.910 1410.670 ;
        RECT 1224.130 1231.090 1225.310 1232.270 ;
        RECT 1225.730 1231.090 1226.910 1232.270 ;
        RECT 1224.130 1229.490 1225.310 1230.670 ;
        RECT 1225.730 1229.490 1226.910 1230.670 ;
        RECT 1224.130 1051.090 1225.310 1052.270 ;
        RECT 1225.730 1051.090 1226.910 1052.270 ;
        RECT 1224.130 1049.490 1225.310 1050.670 ;
        RECT 1225.730 1049.490 1226.910 1050.670 ;
        RECT 1224.130 871.090 1225.310 872.270 ;
        RECT 1225.730 871.090 1226.910 872.270 ;
        RECT 1224.130 869.490 1225.310 870.670 ;
        RECT 1225.730 869.490 1226.910 870.670 ;
        RECT 1224.130 691.090 1225.310 692.270 ;
        RECT 1225.730 691.090 1226.910 692.270 ;
        RECT 1224.130 689.490 1225.310 690.670 ;
        RECT 1225.730 689.490 1226.910 690.670 ;
        RECT 1224.130 511.090 1225.310 512.270 ;
        RECT 1225.730 511.090 1226.910 512.270 ;
        RECT 1224.130 509.490 1225.310 510.670 ;
        RECT 1225.730 509.490 1226.910 510.670 ;
        RECT 1224.130 331.090 1225.310 332.270 ;
        RECT 1225.730 331.090 1226.910 332.270 ;
        RECT 1224.130 329.490 1225.310 330.670 ;
        RECT 1225.730 329.490 1226.910 330.670 ;
        RECT 1224.130 151.090 1225.310 152.270 ;
        RECT 1225.730 151.090 1226.910 152.270 ;
        RECT 1224.130 149.490 1225.310 150.670 ;
        RECT 1225.730 149.490 1226.910 150.670 ;
        RECT 1224.130 -31.710 1225.310 -30.530 ;
        RECT 1225.730 -31.710 1226.910 -30.530 ;
        RECT 1224.130 -33.310 1225.310 -32.130 ;
        RECT 1225.730 -33.310 1226.910 -32.130 ;
        RECT 1404.130 3551.810 1405.310 3552.990 ;
        RECT 1405.730 3551.810 1406.910 3552.990 ;
        RECT 1404.130 3550.210 1405.310 3551.390 ;
        RECT 1405.730 3550.210 1406.910 3551.390 ;
        RECT 1404.130 3391.090 1405.310 3392.270 ;
        RECT 1405.730 3391.090 1406.910 3392.270 ;
        RECT 1404.130 3389.490 1405.310 3390.670 ;
        RECT 1405.730 3389.490 1406.910 3390.670 ;
        RECT 1404.130 3211.090 1405.310 3212.270 ;
        RECT 1405.730 3211.090 1406.910 3212.270 ;
        RECT 1404.130 3209.490 1405.310 3210.670 ;
        RECT 1405.730 3209.490 1406.910 3210.670 ;
        RECT 1404.130 3031.090 1405.310 3032.270 ;
        RECT 1405.730 3031.090 1406.910 3032.270 ;
        RECT 1404.130 3029.490 1405.310 3030.670 ;
        RECT 1405.730 3029.490 1406.910 3030.670 ;
        RECT 1404.130 2851.090 1405.310 2852.270 ;
        RECT 1405.730 2851.090 1406.910 2852.270 ;
        RECT 1404.130 2849.490 1405.310 2850.670 ;
        RECT 1405.730 2849.490 1406.910 2850.670 ;
        RECT 1404.130 2671.090 1405.310 2672.270 ;
        RECT 1405.730 2671.090 1406.910 2672.270 ;
        RECT 1404.130 2669.490 1405.310 2670.670 ;
        RECT 1405.730 2669.490 1406.910 2670.670 ;
        RECT 1404.130 2491.090 1405.310 2492.270 ;
        RECT 1405.730 2491.090 1406.910 2492.270 ;
        RECT 1404.130 2489.490 1405.310 2490.670 ;
        RECT 1405.730 2489.490 1406.910 2490.670 ;
        RECT 1404.130 2311.090 1405.310 2312.270 ;
        RECT 1405.730 2311.090 1406.910 2312.270 ;
        RECT 1404.130 2309.490 1405.310 2310.670 ;
        RECT 1405.730 2309.490 1406.910 2310.670 ;
        RECT 1404.130 2131.090 1405.310 2132.270 ;
        RECT 1405.730 2131.090 1406.910 2132.270 ;
        RECT 1404.130 2129.490 1405.310 2130.670 ;
        RECT 1405.730 2129.490 1406.910 2130.670 ;
        RECT 1404.130 1951.090 1405.310 1952.270 ;
        RECT 1405.730 1951.090 1406.910 1952.270 ;
        RECT 1404.130 1949.490 1405.310 1950.670 ;
        RECT 1405.730 1949.490 1406.910 1950.670 ;
        RECT 1404.130 1771.090 1405.310 1772.270 ;
        RECT 1405.730 1771.090 1406.910 1772.270 ;
        RECT 1404.130 1769.490 1405.310 1770.670 ;
        RECT 1405.730 1769.490 1406.910 1770.670 ;
        RECT 1404.130 1591.090 1405.310 1592.270 ;
        RECT 1405.730 1591.090 1406.910 1592.270 ;
        RECT 1404.130 1589.490 1405.310 1590.670 ;
        RECT 1405.730 1589.490 1406.910 1590.670 ;
        RECT 1404.130 1411.090 1405.310 1412.270 ;
        RECT 1405.730 1411.090 1406.910 1412.270 ;
        RECT 1404.130 1409.490 1405.310 1410.670 ;
        RECT 1405.730 1409.490 1406.910 1410.670 ;
        RECT 1404.130 1231.090 1405.310 1232.270 ;
        RECT 1405.730 1231.090 1406.910 1232.270 ;
        RECT 1404.130 1229.490 1405.310 1230.670 ;
        RECT 1405.730 1229.490 1406.910 1230.670 ;
        RECT 1404.130 1051.090 1405.310 1052.270 ;
        RECT 1405.730 1051.090 1406.910 1052.270 ;
        RECT 1404.130 1049.490 1405.310 1050.670 ;
        RECT 1405.730 1049.490 1406.910 1050.670 ;
        RECT 1404.130 871.090 1405.310 872.270 ;
        RECT 1405.730 871.090 1406.910 872.270 ;
        RECT 1404.130 869.490 1405.310 870.670 ;
        RECT 1405.730 869.490 1406.910 870.670 ;
        RECT 1404.130 691.090 1405.310 692.270 ;
        RECT 1405.730 691.090 1406.910 692.270 ;
        RECT 1404.130 689.490 1405.310 690.670 ;
        RECT 1405.730 689.490 1406.910 690.670 ;
        RECT 1404.130 511.090 1405.310 512.270 ;
        RECT 1405.730 511.090 1406.910 512.270 ;
        RECT 1404.130 509.490 1405.310 510.670 ;
        RECT 1405.730 509.490 1406.910 510.670 ;
        RECT 1404.130 331.090 1405.310 332.270 ;
        RECT 1405.730 331.090 1406.910 332.270 ;
        RECT 1404.130 329.490 1405.310 330.670 ;
        RECT 1405.730 329.490 1406.910 330.670 ;
        RECT 1404.130 151.090 1405.310 152.270 ;
        RECT 1405.730 151.090 1406.910 152.270 ;
        RECT 1404.130 149.490 1405.310 150.670 ;
        RECT 1405.730 149.490 1406.910 150.670 ;
        RECT 1404.130 -31.710 1405.310 -30.530 ;
        RECT 1405.730 -31.710 1406.910 -30.530 ;
        RECT 1404.130 -33.310 1405.310 -32.130 ;
        RECT 1405.730 -33.310 1406.910 -32.130 ;
        RECT 1584.130 3551.810 1585.310 3552.990 ;
        RECT 1585.730 3551.810 1586.910 3552.990 ;
        RECT 1584.130 3550.210 1585.310 3551.390 ;
        RECT 1585.730 3550.210 1586.910 3551.390 ;
        RECT 1584.130 3391.090 1585.310 3392.270 ;
        RECT 1585.730 3391.090 1586.910 3392.270 ;
        RECT 1584.130 3389.490 1585.310 3390.670 ;
        RECT 1585.730 3389.490 1586.910 3390.670 ;
        RECT 1584.130 3211.090 1585.310 3212.270 ;
        RECT 1585.730 3211.090 1586.910 3212.270 ;
        RECT 1584.130 3209.490 1585.310 3210.670 ;
        RECT 1585.730 3209.490 1586.910 3210.670 ;
        RECT 1584.130 3031.090 1585.310 3032.270 ;
        RECT 1585.730 3031.090 1586.910 3032.270 ;
        RECT 1584.130 3029.490 1585.310 3030.670 ;
        RECT 1585.730 3029.490 1586.910 3030.670 ;
        RECT 1584.130 2851.090 1585.310 2852.270 ;
        RECT 1585.730 2851.090 1586.910 2852.270 ;
        RECT 1584.130 2849.490 1585.310 2850.670 ;
        RECT 1585.730 2849.490 1586.910 2850.670 ;
        RECT 1584.130 2671.090 1585.310 2672.270 ;
        RECT 1585.730 2671.090 1586.910 2672.270 ;
        RECT 1584.130 2669.490 1585.310 2670.670 ;
        RECT 1585.730 2669.490 1586.910 2670.670 ;
        RECT 1584.130 2491.090 1585.310 2492.270 ;
        RECT 1585.730 2491.090 1586.910 2492.270 ;
        RECT 1584.130 2489.490 1585.310 2490.670 ;
        RECT 1585.730 2489.490 1586.910 2490.670 ;
        RECT 1584.130 2311.090 1585.310 2312.270 ;
        RECT 1585.730 2311.090 1586.910 2312.270 ;
        RECT 1584.130 2309.490 1585.310 2310.670 ;
        RECT 1585.730 2309.490 1586.910 2310.670 ;
        RECT 1584.130 2131.090 1585.310 2132.270 ;
        RECT 1585.730 2131.090 1586.910 2132.270 ;
        RECT 1584.130 2129.490 1585.310 2130.670 ;
        RECT 1585.730 2129.490 1586.910 2130.670 ;
        RECT 1584.130 1951.090 1585.310 1952.270 ;
        RECT 1585.730 1951.090 1586.910 1952.270 ;
        RECT 1584.130 1949.490 1585.310 1950.670 ;
        RECT 1585.730 1949.490 1586.910 1950.670 ;
        RECT 1584.130 1771.090 1585.310 1772.270 ;
        RECT 1585.730 1771.090 1586.910 1772.270 ;
        RECT 1584.130 1769.490 1585.310 1770.670 ;
        RECT 1585.730 1769.490 1586.910 1770.670 ;
        RECT 1584.130 1591.090 1585.310 1592.270 ;
        RECT 1585.730 1591.090 1586.910 1592.270 ;
        RECT 1584.130 1589.490 1585.310 1590.670 ;
        RECT 1585.730 1589.490 1586.910 1590.670 ;
        RECT 1584.130 1411.090 1585.310 1412.270 ;
        RECT 1585.730 1411.090 1586.910 1412.270 ;
        RECT 1584.130 1409.490 1585.310 1410.670 ;
        RECT 1585.730 1409.490 1586.910 1410.670 ;
        RECT 1584.130 1231.090 1585.310 1232.270 ;
        RECT 1585.730 1231.090 1586.910 1232.270 ;
        RECT 1584.130 1229.490 1585.310 1230.670 ;
        RECT 1585.730 1229.490 1586.910 1230.670 ;
        RECT 1584.130 1051.090 1585.310 1052.270 ;
        RECT 1585.730 1051.090 1586.910 1052.270 ;
        RECT 1584.130 1049.490 1585.310 1050.670 ;
        RECT 1585.730 1049.490 1586.910 1050.670 ;
        RECT 1584.130 871.090 1585.310 872.270 ;
        RECT 1585.730 871.090 1586.910 872.270 ;
        RECT 1584.130 869.490 1585.310 870.670 ;
        RECT 1585.730 869.490 1586.910 870.670 ;
        RECT 1584.130 691.090 1585.310 692.270 ;
        RECT 1585.730 691.090 1586.910 692.270 ;
        RECT 1584.130 689.490 1585.310 690.670 ;
        RECT 1585.730 689.490 1586.910 690.670 ;
        RECT 1584.130 511.090 1585.310 512.270 ;
        RECT 1585.730 511.090 1586.910 512.270 ;
        RECT 1584.130 509.490 1585.310 510.670 ;
        RECT 1585.730 509.490 1586.910 510.670 ;
        RECT 1584.130 331.090 1585.310 332.270 ;
        RECT 1585.730 331.090 1586.910 332.270 ;
        RECT 1584.130 329.490 1585.310 330.670 ;
        RECT 1585.730 329.490 1586.910 330.670 ;
        RECT 1584.130 151.090 1585.310 152.270 ;
        RECT 1585.730 151.090 1586.910 152.270 ;
        RECT 1584.130 149.490 1585.310 150.670 ;
        RECT 1585.730 149.490 1586.910 150.670 ;
        RECT 1584.130 -31.710 1585.310 -30.530 ;
        RECT 1585.730 -31.710 1586.910 -30.530 ;
        RECT 1584.130 -33.310 1585.310 -32.130 ;
        RECT 1585.730 -33.310 1586.910 -32.130 ;
        RECT 1764.130 3551.810 1765.310 3552.990 ;
        RECT 1765.730 3551.810 1766.910 3552.990 ;
        RECT 1764.130 3550.210 1765.310 3551.390 ;
        RECT 1765.730 3550.210 1766.910 3551.390 ;
        RECT 1764.130 3391.090 1765.310 3392.270 ;
        RECT 1765.730 3391.090 1766.910 3392.270 ;
        RECT 1764.130 3389.490 1765.310 3390.670 ;
        RECT 1765.730 3389.490 1766.910 3390.670 ;
        RECT 1764.130 3211.090 1765.310 3212.270 ;
        RECT 1765.730 3211.090 1766.910 3212.270 ;
        RECT 1764.130 3209.490 1765.310 3210.670 ;
        RECT 1765.730 3209.490 1766.910 3210.670 ;
        RECT 1764.130 3031.090 1765.310 3032.270 ;
        RECT 1765.730 3031.090 1766.910 3032.270 ;
        RECT 1764.130 3029.490 1765.310 3030.670 ;
        RECT 1765.730 3029.490 1766.910 3030.670 ;
        RECT 1764.130 2851.090 1765.310 2852.270 ;
        RECT 1765.730 2851.090 1766.910 2852.270 ;
        RECT 1764.130 2849.490 1765.310 2850.670 ;
        RECT 1765.730 2849.490 1766.910 2850.670 ;
        RECT 1764.130 2671.090 1765.310 2672.270 ;
        RECT 1765.730 2671.090 1766.910 2672.270 ;
        RECT 1764.130 2669.490 1765.310 2670.670 ;
        RECT 1765.730 2669.490 1766.910 2670.670 ;
        RECT 1764.130 2491.090 1765.310 2492.270 ;
        RECT 1765.730 2491.090 1766.910 2492.270 ;
        RECT 1764.130 2489.490 1765.310 2490.670 ;
        RECT 1765.730 2489.490 1766.910 2490.670 ;
        RECT 1764.130 2311.090 1765.310 2312.270 ;
        RECT 1765.730 2311.090 1766.910 2312.270 ;
        RECT 1764.130 2309.490 1765.310 2310.670 ;
        RECT 1765.730 2309.490 1766.910 2310.670 ;
        RECT 1764.130 2131.090 1765.310 2132.270 ;
        RECT 1765.730 2131.090 1766.910 2132.270 ;
        RECT 1764.130 2129.490 1765.310 2130.670 ;
        RECT 1765.730 2129.490 1766.910 2130.670 ;
        RECT 1764.130 1951.090 1765.310 1952.270 ;
        RECT 1765.730 1951.090 1766.910 1952.270 ;
        RECT 1764.130 1949.490 1765.310 1950.670 ;
        RECT 1765.730 1949.490 1766.910 1950.670 ;
        RECT 1764.130 1771.090 1765.310 1772.270 ;
        RECT 1765.730 1771.090 1766.910 1772.270 ;
        RECT 1764.130 1769.490 1765.310 1770.670 ;
        RECT 1765.730 1769.490 1766.910 1770.670 ;
        RECT 1764.130 1591.090 1765.310 1592.270 ;
        RECT 1765.730 1591.090 1766.910 1592.270 ;
        RECT 1764.130 1589.490 1765.310 1590.670 ;
        RECT 1765.730 1589.490 1766.910 1590.670 ;
        RECT 1764.130 1411.090 1765.310 1412.270 ;
        RECT 1765.730 1411.090 1766.910 1412.270 ;
        RECT 1764.130 1409.490 1765.310 1410.670 ;
        RECT 1765.730 1409.490 1766.910 1410.670 ;
        RECT 1764.130 1231.090 1765.310 1232.270 ;
        RECT 1765.730 1231.090 1766.910 1232.270 ;
        RECT 1764.130 1229.490 1765.310 1230.670 ;
        RECT 1765.730 1229.490 1766.910 1230.670 ;
        RECT 1764.130 1051.090 1765.310 1052.270 ;
        RECT 1765.730 1051.090 1766.910 1052.270 ;
        RECT 1764.130 1049.490 1765.310 1050.670 ;
        RECT 1765.730 1049.490 1766.910 1050.670 ;
        RECT 1764.130 871.090 1765.310 872.270 ;
        RECT 1765.730 871.090 1766.910 872.270 ;
        RECT 1764.130 869.490 1765.310 870.670 ;
        RECT 1765.730 869.490 1766.910 870.670 ;
        RECT 1764.130 691.090 1765.310 692.270 ;
        RECT 1765.730 691.090 1766.910 692.270 ;
        RECT 1764.130 689.490 1765.310 690.670 ;
        RECT 1765.730 689.490 1766.910 690.670 ;
        RECT 1764.130 511.090 1765.310 512.270 ;
        RECT 1765.730 511.090 1766.910 512.270 ;
        RECT 1764.130 509.490 1765.310 510.670 ;
        RECT 1765.730 509.490 1766.910 510.670 ;
        RECT 1764.130 331.090 1765.310 332.270 ;
        RECT 1765.730 331.090 1766.910 332.270 ;
        RECT 1764.130 329.490 1765.310 330.670 ;
        RECT 1765.730 329.490 1766.910 330.670 ;
        RECT 1764.130 151.090 1765.310 152.270 ;
        RECT 1765.730 151.090 1766.910 152.270 ;
        RECT 1764.130 149.490 1765.310 150.670 ;
        RECT 1765.730 149.490 1766.910 150.670 ;
        RECT 1764.130 -31.710 1765.310 -30.530 ;
        RECT 1765.730 -31.710 1766.910 -30.530 ;
        RECT 1764.130 -33.310 1765.310 -32.130 ;
        RECT 1765.730 -33.310 1766.910 -32.130 ;
        RECT 1944.130 3551.810 1945.310 3552.990 ;
        RECT 1945.730 3551.810 1946.910 3552.990 ;
        RECT 1944.130 3550.210 1945.310 3551.390 ;
        RECT 1945.730 3550.210 1946.910 3551.390 ;
        RECT 1944.130 3391.090 1945.310 3392.270 ;
        RECT 1945.730 3391.090 1946.910 3392.270 ;
        RECT 1944.130 3389.490 1945.310 3390.670 ;
        RECT 1945.730 3389.490 1946.910 3390.670 ;
        RECT 1944.130 3211.090 1945.310 3212.270 ;
        RECT 1945.730 3211.090 1946.910 3212.270 ;
        RECT 1944.130 3209.490 1945.310 3210.670 ;
        RECT 1945.730 3209.490 1946.910 3210.670 ;
        RECT 1944.130 3031.090 1945.310 3032.270 ;
        RECT 1945.730 3031.090 1946.910 3032.270 ;
        RECT 1944.130 3029.490 1945.310 3030.670 ;
        RECT 1945.730 3029.490 1946.910 3030.670 ;
        RECT 1944.130 2851.090 1945.310 2852.270 ;
        RECT 1945.730 2851.090 1946.910 2852.270 ;
        RECT 1944.130 2849.490 1945.310 2850.670 ;
        RECT 1945.730 2849.490 1946.910 2850.670 ;
        RECT 1944.130 2671.090 1945.310 2672.270 ;
        RECT 1945.730 2671.090 1946.910 2672.270 ;
        RECT 1944.130 2669.490 1945.310 2670.670 ;
        RECT 1945.730 2669.490 1946.910 2670.670 ;
        RECT 1944.130 2491.090 1945.310 2492.270 ;
        RECT 1945.730 2491.090 1946.910 2492.270 ;
        RECT 1944.130 2489.490 1945.310 2490.670 ;
        RECT 1945.730 2489.490 1946.910 2490.670 ;
        RECT 1944.130 2311.090 1945.310 2312.270 ;
        RECT 1945.730 2311.090 1946.910 2312.270 ;
        RECT 1944.130 2309.490 1945.310 2310.670 ;
        RECT 1945.730 2309.490 1946.910 2310.670 ;
        RECT 1944.130 2131.090 1945.310 2132.270 ;
        RECT 1945.730 2131.090 1946.910 2132.270 ;
        RECT 1944.130 2129.490 1945.310 2130.670 ;
        RECT 1945.730 2129.490 1946.910 2130.670 ;
        RECT 1944.130 1951.090 1945.310 1952.270 ;
        RECT 1945.730 1951.090 1946.910 1952.270 ;
        RECT 1944.130 1949.490 1945.310 1950.670 ;
        RECT 1945.730 1949.490 1946.910 1950.670 ;
        RECT 1944.130 1771.090 1945.310 1772.270 ;
        RECT 1945.730 1771.090 1946.910 1772.270 ;
        RECT 1944.130 1769.490 1945.310 1770.670 ;
        RECT 1945.730 1769.490 1946.910 1770.670 ;
        RECT 1944.130 1591.090 1945.310 1592.270 ;
        RECT 1945.730 1591.090 1946.910 1592.270 ;
        RECT 1944.130 1589.490 1945.310 1590.670 ;
        RECT 1945.730 1589.490 1946.910 1590.670 ;
        RECT 1944.130 1411.090 1945.310 1412.270 ;
        RECT 1945.730 1411.090 1946.910 1412.270 ;
        RECT 1944.130 1409.490 1945.310 1410.670 ;
        RECT 1945.730 1409.490 1946.910 1410.670 ;
        RECT 1944.130 1231.090 1945.310 1232.270 ;
        RECT 1945.730 1231.090 1946.910 1232.270 ;
        RECT 1944.130 1229.490 1945.310 1230.670 ;
        RECT 1945.730 1229.490 1946.910 1230.670 ;
        RECT 1944.130 1051.090 1945.310 1052.270 ;
        RECT 1945.730 1051.090 1946.910 1052.270 ;
        RECT 1944.130 1049.490 1945.310 1050.670 ;
        RECT 1945.730 1049.490 1946.910 1050.670 ;
        RECT 1944.130 871.090 1945.310 872.270 ;
        RECT 1945.730 871.090 1946.910 872.270 ;
        RECT 1944.130 869.490 1945.310 870.670 ;
        RECT 1945.730 869.490 1946.910 870.670 ;
        RECT 1944.130 691.090 1945.310 692.270 ;
        RECT 1945.730 691.090 1946.910 692.270 ;
        RECT 1944.130 689.490 1945.310 690.670 ;
        RECT 1945.730 689.490 1946.910 690.670 ;
        RECT 1944.130 511.090 1945.310 512.270 ;
        RECT 1945.730 511.090 1946.910 512.270 ;
        RECT 1944.130 509.490 1945.310 510.670 ;
        RECT 1945.730 509.490 1946.910 510.670 ;
        RECT 1944.130 331.090 1945.310 332.270 ;
        RECT 1945.730 331.090 1946.910 332.270 ;
        RECT 1944.130 329.490 1945.310 330.670 ;
        RECT 1945.730 329.490 1946.910 330.670 ;
        RECT 1944.130 151.090 1945.310 152.270 ;
        RECT 1945.730 151.090 1946.910 152.270 ;
        RECT 1944.130 149.490 1945.310 150.670 ;
        RECT 1945.730 149.490 1946.910 150.670 ;
        RECT 1944.130 -31.710 1945.310 -30.530 ;
        RECT 1945.730 -31.710 1946.910 -30.530 ;
        RECT 1944.130 -33.310 1945.310 -32.130 ;
        RECT 1945.730 -33.310 1946.910 -32.130 ;
        RECT 2124.130 3551.810 2125.310 3552.990 ;
        RECT 2125.730 3551.810 2126.910 3552.990 ;
        RECT 2124.130 3550.210 2125.310 3551.390 ;
        RECT 2125.730 3550.210 2126.910 3551.390 ;
        RECT 2124.130 3391.090 2125.310 3392.270 ;
        RECT 2125.730 3391.090 2126.910 3392.270 ;
        RECT 2124.130 3389.490 2125.310 3390.670 ;
        RECT 2125.730 3389.490 2126.910 3390.670 ;
        RECT 2124.130 3211.090 2125.310 3212.270 ;
        RECT 2125.730 3211.090 2126.910 3212.270 ;
        RECT 2124.130 3209.490 2125.310 3210.670 ;
        RECT 2125.730 3209.490 2126.910 3210.670 ;
        RECT 2124.130 3031.090 2125.310 3032.270 ;
        RECT 2125.730 3031.090 2126.910 3032.270 ;
        RECT 2124.130 3029.490 2125.310 3030.670 ;
        RECT 2125.730 3029.490 2126.910 3030.670 ;
        RECT 2124.130 2851.090 2125.310 2852.270 ;
        RECT 2125.730 2851.090 2126.910 2852.270 ;
        RECT 2124.130 2849.490 2125.310 2850.670 ;
        RECT 2125.730 2849.490 2126.910 2850.670 ;
        RECT 2124.130 2671.090 2125.310 2672.270 ;
        RECT 2125.730 2671.090 2126.910 2672.270 ;
        RECT 2124.130 2669.490 2125.310 2670.670 ;
        RECT 2125.730 2669.490 2126.910 2670.670 ;
        RECT 2124.130 2491.090 2125.310 2492.270 ;
        RECT 2125.730 2491.090 2126.910 2492.270 ;
        RECT 2124.130 2489.490 2125.310 2490.670 ;
        RECT 2125.730 2489.490 2126.910 2490.670 ;
        RECT 2124.130 2311.090 2125.310 2312.270 ;
        RECT 2125.730 2311.090 2126.910 2312.270 ;
        RECT 2124.130 2309.490 2125.310 2310.670 ;
        RECT 2125.730 2309.490 2126.910 2310.670 ;
        RECT 2124.130 2131.090 2125.310 2132.270 ;
        RECT 2125.730 2131.090 2126.910 2132.270 ;
        RECT 2124.130 2129.490 2125.310 2130.670 ;
        RECT 2125.730 2129.490 2126.910 2130.670 ;
        RECT 2124.130 1951.090 2125.310 1952.270 ;
        RECT 2125.730 1951.090 2126.910 1952.270 ;
        RECT 2124.130 1949.490 2125.310 1950.670 ;
        RECT 2125.730 1949.490 2126.910 1950.670 ;
        RECT 2124.130 1771.090 2125.310 1772.270 ;
        RECT 2125.730 1771.090 2126.910 1772.270 ;
        RECT 2124.130 1769.490 2125.310 1770.670 ;
        RECT 2125.730 1769.490 2126.910 1770.670 ;
        RECT 2124.130 1591.090 2125.310 1592.270 ;
        RECT 2125.730 1591.090 2126.910 1592.270 ;
        RECT 2124.130 1589.490 2125.310 1590.670 ;
        RECT 2125.730 1589.490 2126.910 1590.670 ;
        RECT 2124.130 1411.090 2125.310 1412.270 ;
        RECT 2125.730 1411.090 2126.910 1412.270 ;
        RECT 2124.130 1409.490 2125.310 1410.670 ;
        RECT 2125.730 1409.490 2126.910 1410.670 ;
        RECT 2124.130 1231.090 2125.310 1232.270 ;
        RECT 2125.730 1231.090 2126.910 1232.270 ;
        RECT 2124.130 1229.490 2125.310 1230.670 ;
        RECT 2125.730 1229.490 2126.910 1230.670 ;
        RECT 2124.130 1051.090 2125.310 1052.270 ;
        RECT 2125.730 1051.090 2126.910 1052.270 ;
        RECT 2124.130 1049.490 2125.310 1050.670 ;
        RECT 2125.730 1049.490 2126.910 1050.670 ;
        RECT 2124.130 871.090 2125.310 872.270 ;
        RECT 2125.730 871.090 2126.910 872.270 ;
        RECT 2124.130 869.490 2125.310 870.670 ;
        RECT 2125.730 869.490 2126.910 870.670 ;
        RECT 2124.130 691.090 2125.310 692.270 ;
        RECT 2125.730 691.090 2126.910 692.270 ;
        RECT 2124.130 689.490 2125.310 690.670 ;
        RECT 2125.730 689.490 2126.910 690.670 ;
        RECT 2124.130 511.090 2125.310 512.270 ;
        RECT 2125.730 511.090 2126.910 512.270 ;
        RECT 2124.130 509.490 2125.310 510.670 ;
        RECT 2125.730 509.490 2126.910 510.670 ;
        RECT 2124.130 331.090 2125.310 332.270 ;
        RECT 2125.730 331.090 2126.910 332.270 ;
        RECT 2124.130 329.490 2125.310 330.670 ;
        RECT 2125.730 329.490 2126.910 330.670 ;
        RECT 2124.130 151.090 2125.310 152.270 ;
        RECT 2125.730 151.090 2126.910 152.270 ;
        RECT 2124.130 149.490 2125.310 150.670 ;
        RECT 2125.730 149.490 2126.910 150.670 ;
        RECT 2124.130 -31.710 2125.310 -30.530 ;
        RECT 2125.730 -31.710 2126.910 -30.530 ;
        RECT 2124.130 -33.310 2125.310 -32.130 ;
        RECT 2125.730 -33.310 2126.910 -32.130 ;
        RECT 2304.130 3551.810 2305.310 3552.990 ;
        RECT 2305.730 3551.810 2306.910 3552.990 ;
        RECT 2304.130 3550.210 2305.310 3551.390 ;
        RECT 2305.730 3550.210 2306.910 3551.390 ;
        RECT 2304.130 3391.090 2305.310 3392.270 ;
        RECT 2305.730 3391.090 2306.910 3392.270 ;
        RECT 2304.130 3389.490 2305.310 3390.670 ;
        RECT 2305.730 3389.490 2306.910 3390.670 ;
        RECT 2304.130 3211.090 2305.310 3212.270 ;
        RECT 2305.730 3211.090 2306.910 3212.270 ;
        RECT 2304.130 3209.490 2305.310 3210.670 ;
        RECT 2305.730 3209.490 2306.910 3210.670 ;
        RECT 2304.130 3031.090 2305.310 3032.270 ;
        RECT 2305.730 3031.090 2306.910 3032.270 ;
        RECT 2304.130 3029.490 2305.310 3030.670 ;
        RECT 2305.730 3029.490 2306.910 3030.670 ;
        RECT 2304.130 2851.090 2305.310 2852.270 ;
        RECT 2305.730 2851.090 2306.910 2852.270 ;
        RECT 2304.130 2849.490 2305.310 2850.670 ;
        RECT 2305.730 2849.490 2306.910 2850.670 ;
        RECT 2304.130 2671.090 2305.310 2672.270 ;
        RECT 2305.730 2671.090 2306.910 2672.270 ;
        RECT 2304.130 2669.490 2305.310 2670.670 ;
        RECT 2305.730 2669.490 2306.910 2670.670 ;
        RECT 2304.130 2491.090 2305.310 2492.270 ;
        RECT 2305.730 2491.090 2306.910 2492.270 ;
        RECT 2304.130 2489.490 2305.310 2490.670 ;
        RECT 2305.730 2489.490 2306.910 2490.670 ;
        RECT 2304.130 2311.090 2305.310 2312.270 ;
        RECT 2305.730 2311.090 2306.910 2312.270 ;
        RECT 2304.130 2309.490 2305.310 2310.670 ;
        RECT 2305.730 2309.490 2306.910 2310.670 ;
        RECT 2304.130 2131.090 2305.310 2132.270 ;
        RECT 2305.730 2131.090 2306.910 2132.270 ;
        RECT 2304.130 2129.490 2305.310 2130.670 ;
        RECT 2305.730 2129.490 2306.910 2130.670 ;
        RECT 2304.130 1951.090 2305.310 1952.270 ;
        RECT 2305.730 1951.090 2306.910 1952.270 ;
        RECT 2304.130 1949.490 2305.310 1950.670 ;
        RECT 2305.730 1949.490 2306.910 1950.670 ;
        RECT 2304.130 1771.090 2305.310 1772.270 ;
        RECT 2305.730 1771.090 2306.910 1772.270 ;
        RECT 2304.130 1769.490 2305.310 1770.670 ;
        RECT 2305.730 1769.490 2306.910 1770.670 ;
        RECT 2304.130 1591.090 2305.310 1592.270 ;
        RECT 2305.730 1591.090 2306.910 1592.270 ;
        RECT 2304.130 1589.490 2305.310 1590.670 ;
        RECT 2305.730 1589.490 2306.910 1590.670 ;
        RECT 2304.130 1411.090 2305.310 1412.270 ;
        RECT 2305.730 1411.090 2306.910 1412.270 ;
        RECT 2304.130 1409.490 2305.310 1410.670 ;
        RECT 2305.730 1409.490 2306.910 1410.670 ;
        RECT 2304.130 1231.090 2305.310 1232.270 ;
        RECT 2305.730 1231.090 2306.910 1232.270 ;
        RECT 2304.130 1229.490 2305.310 1230.670 ;
        RECT 2305.730 1229.490 2306.910 1230.670 ;
        RECT 2304.130 1051.090 2305.310 1052.270 ;
        RECT 2305.730 1051.090 2306.910 1052.270 ;
        RECT 2304.130 1049.490 2305.310 1050.670 ;
        RECT 2305.730 1049.490 2306.910 1050.670 ;
        RECT 2304.130 871.090 2305.310 872.270 ;
        RECT 2305.730 871.090 2306.910 872.270 ;
        RECT 2304.130 869.490 2305.310 870.670 ;
        RECT 2305.730 869.490 2306.910 870.670 ;
        RECT 2304.130 691.090 2305.310 692.270 ;
        RECT 2305.730 691.090 2306.910 692.270 ;
        RECT 2304.130 689.490 2305.310 690.670 ;
        RECT 2305.730 689.490 2306.910 690.670 ;
        RECT 2304.130 511.090 2305.310 512.270 ;
        RECT 2305.730 511.090 2306.910 512.270 ;
        RECT 2304.130 509.490 2305.310 510.670 ;
        RECT 2305.730 509.490 2306.910 510.670 ;
        RECT 2304.130 331.090 2305.310 332.270 ;
        RECT 2305.730 331.090 2306.910 332.270 ;
        RECT 2304.130 329.490 2305.310 330.670 ;
        RECT 2305.730 329.490 2306.910 330.670 ;
        RECT 2304.130 151.090 2305.310 152.270 ;
        RECT 2305.730 151.090 2306.910 152.270 ;
        RECT 2304.130 149.490 2305.310 150.670 ;
        RECT 2305.730 149.490 2306.910 150.670 ;
        RECT 2304.130 -31.710 2305.310 -30.530 ;
        RECT 2305.730 -31.710 2306.910 -30.530 ;
        RECT 2304.130 -33.310 2305.310 -32.130 ;
        RECT 2305.730 -33.310 2306.910 -32.130 ;
        RECT 2484.130 3551.810 2485.310 3552.990 ;
        RECT 2485.730 3551.810 2486.910 3552.990 ;
        RECT 2484.130 3550.210 2485.310 3551.390 ;
        RECT 2485.730 3550.210 2486.910 3551.390 ;
        RECT 2484.130 3391.090 2485.310 3392.270 ;
        RECT 2485.730 3391.090 2486.910 3392.270 ;
        RECT 2484.130 3389.490 2485.310 3390.670 ;
        RECT 2485.730 3389.490 2486.910 3390.670 ;
        RECT 2484.130 3211.090 2485.310 3212.270 ;
        RECT 2485.730 3211.090 2486.910 3212.270 ;
        RECT 2484.130 3209.490 2485.310 3210.670 ;
        RECT 2485.730 3209.490 2486.910 3210.670 ;
        RECT 2484.130 3031.090 2485.310 3032.270 ;
        RECT 2485.730 3031.090 2486.910 3032.270 ;
        RECT 2484.130 3029.490 2485.310 3030.670 ;
        RECT 2485.730 3029.490 2486.910 3030.670 ;
        RECT 2484.130 2851.090 2485.310 2852.270 ;
        RECT 2485.730 2851.090 2486.910 2852.270 ;
        RECT 2484.130 2849.490 2485.310 2850.670 ;
        RECT 2485.730 2849.490 2486.910 2850.670 ;
        RECT 2484.130 2671.090 2485.310 2672.270 ;
        RECT 2485.730 2671.090 2486.910 2672.270 ;
        RECT 2484.130 2669.490 2485.310 2670.670 ;
        RECT 2485.730 2669.490 2486.910 2670.670 ;
        RECT 2484.130 2491.090 2485.310 2492.270 ;
        RECT 2485.730 2491.090 2486.910 2492.270 ;
        RECT 2484.130 2489.490 2485.310 2490.670 ;
        RECT 2485.730 2489.490 2486.910 2490.670 ;
        RECT 2484.130 2311.090 2485.310 2312.270 ;
        RECT 2485.730 2311.090 2486.910 2312.270 ;
        RECT 2484.130 2309.490 2485.310 2310.670 ;
        RECT 2485.730 2309.490 2486.910 2310.670 ;
        RECT 2484.130 2131.090 2485.310 2132.270 ;
        RECT 2485.730 2131.090 2486.910 2132.270 ;
        RECT 2484.130 2129.490 2485.310 2130.670 ;
        RECT 2485.730 2129.490 2486.910 2130.670 ;
        RECT 2484.130 1951.090 2485.310 1952.270 ;
        RECT 2485.730 1951.090 2486.910 1952.270 ;
        RECT 2484.130 1949.490 2485.310 1950.670 ;
        RECT 2485.730 1949.490 2486.910 1950.670 ;
        RECT 2484.130 1771.090 2485.310 1772.270 ;
        RECT 2485.730 1771.090 2486.910 1772.270 ;
        RECT 2484.130 1769.490 2485.310 1770.670 ;
        RECT 2485.730 1769.490 2486.910 1770.670 ;
        RECT 2484.130 1591.090 2485.310 1592.270 ;
        RECT 2485.730 1591.090 2486.910 1592.270 ;
        RECT 2484.130 1589.490 2485.310 1590.670 ;
        RECT 2485.730 1589.490 2486.910 1590.670 ;
        RECT 2484.130 1411.090 2485.310 1412.270 ;
        RECT 2485.730 1411.090 2486.910 1412.270 ;
        RECT 2484.130 1409.490 2485.310 1410.670 ;
        RECT 2485.730 1409.490 2486.910 1410.670 ;
        RECT 2484.130 1231.090 2485.310 1232.270 ;
        RECT 2485.730 1231.090 2486.910 1232.270 ;
        RECT 2484.130 1229.490 2485.310 1230.670 ;
        RECT 2485.730 1229.490 2486.910 1230.670 ;
        RECT 2484.130 1051.090 2485.310 1052.270 ;
        RECT 2485.730 1051.090 2486.910 1052.270 ;
        RECT 2484.130 1049.490 2485.310 1050.670 ;
        RECT 2485.730 1049.490 2486.910 1050.670 ;
        RECT 2484.130 871.090 2485.310 872.270 ;
        RECT 2485.730 871.090 2486.910 872.270 ;
        RECT 2484.130 869.490 2485.310 870.670 ;
        RECT 2485.730 869.490 2486.910 870.670 ;
        RECT 2484.130 691.090 2485.310 692.270 ;
        RECT 2485.730 691.090 2486.910 692.270 ;
        RECT 2484.130 689.490 2485.310 690.670 ;
        RECT 2485.730 689.490 2486.910 690.670 ;
        RECT 2484.130 511.090 2485.310 512.270 ;
        RECT 2485.730 511.090 2486.910 512.270 ;
        RECT 2484.130 509.490 2485.310 510.670 ;
        RECT 2485.730 509.490 2486.910 510.670 ;
        RECT 2484.130 331.090 2485.310 332.270 ;
        RECT 2485.730 331.090 2486.910 332.270 ;
        RECT 2484.130 329.490 2485.310 330.670 ;
        RECT 2485.730 329.490 2486.910 330.670 ;
        RECT 2484.130 151.090 2485.310 152.270 ;
        RECT 2485.730 151.090 2486.910 152.270 ;
        RECT 2484.130 149.490 2485.310 150.670 ;
        RECT 2485.730 149.490 2486.910 150.670 ;
        RECT 2484.130 -31.710 2485.310 -30.530 ;
        RECT 2485.730 -31.710 2486.910 -30.530 ;
        RECT 2484.130 -33.310 2485.310 -32.130 ;
        RECT 2485.730 -33.310 2486.910 -32.130 ;
        RECT 2664.130 3551.810 2665.310 3552.990 ;
        RECT 2665.730 3551.810 2666.910 3552.990 ;
        RECT 2664.130 3550.210 2665.310 3551.390 ;
        RECT 2665.730 3550.210 2666.910 3551.390 ;
        RECT 2664.130 3391.090 2665.310 3392.270 ;
        RECT 2665.730 3391.090 2666.910 3392.270 ;
        RECT 2664.130 3389.490 2665.310 3390.670 ;
        RECT 2665.730 3389.490 2666.910 3390.670 ;
        RECT 2664.130 3211.090 2665.310 3212.270 ;
        RECT 2665.730 3211.090 2666.910 3212.270 ;
        RECT 2664.130 3209.490 2665.310 3210.670 ;
        RECT 2665.730 3209.490 2666.910 3210.670 ;
        RECT 2664.130 3031.090 2665.310 3032.270 ;
        RECT 2665.730 3031.090 2666.910 3032.270 ;
        RECT 2664.130 3029.490 2665.310 3030.670 ;
        RECT 2665.730 3029.490 2666.910 3030.670 ;
        RECT 2664.130 2851.090 2665.310 2852.270 ;
        RECT 2665.730 2851.090 2666.910 2852.270 ;
        RECT 2664.130 2849.490 2665.310 2850.670 ;
        RECT 2665.730 2849.490 2666.910 2850.670 ;
        RECT 2664.130 2671.090 2665.310 2672.270 ;
        RECT 2665.730 2671.090 2666.910 2672.270 ;
        RECT 2664.130 2669.490 2665.310 2670.670 ;
        RECT 2665.730 2669.490 2666.910 2670.670 ;
        RECT 2664.130 2491.090 2665.310 2492.270 ;
        RECT 2665.730 2491.090 2666.910 2492.270 ;
        RECT 2664.130 2489.490 2665.310 2490.670 ;
        RECT 2665.730 2489.490 2666.910 2490.670 ;
        RECT 2664.130 2311.090 2665.310 2312.270 ;
        RECT 2665.730 2311.090 2666.910 2312.270 ;
        RECT 2664.130 2309.490 2665.310 2310.670 ;
        RECT 2665.730 2309.490 2666.910 2310.670 ;
        RECT 2664.130 2131.090 2665.310 2132.270 ;
        RECT 2665.730 2131.090 2666.910 2132.270 ;
        RECT 2664.130 2129.490 2665.310 2130.670 ;
        RECT 2665.730 2129.490 2666.910 2130.670 ;
        RECT 2664.130 1951.090 2665.310 1952.270 ;
        RECT 2665.730 1951.090 2666.910 1952.270 ;
        RECT 2664.130 1949.490 2665.310 1950.670 ;
        RECT 2665.730 1949.490 2666.910 1950.670 ;
        RECT 2664.130 1771.090 2665.310 1772.270 ;
        RECT 2665.730 1771.090 2666.910 1772.270 ;
        RECT 2664.130 1769.490 2665.310 1770.670 ;
        RECT 2665.730 1769.490 2666.910 1770.670 ;
        RECT 2664.130 1591.090 2665.310 1592.270 ;
        RECT 2665.730 1591.090 2666.910 1592.270 ;
        RECT 2664.130 1589.490 2665.310 1590.670 ;
        RECT 2665.730 1589.490 2666.910 1590.670 ;
        RECT 2664.130 1411.090 2665.310 1412.270 ;
        RECT 2665.730 1411.090 2666.910 1412.270 ;
        RECT 2664.130 1409.490 2665.310 1410.670 ;
        RECT 2665.730 1409.490 2666.910 1410.670 ;
        RECT 2664.130 1231.090 2665.310 1232.270 ;
        RECT 2665.730 1231.090 2666.910 1232.270 ;
        RECT 2664.130 1229.490 2665.310 1230.670 ;
        RECT 2665.730 1229.490 2666.910 1230.670 ;
        RECT 2664.130 1051.090 2665.310 1052.270 ;
        RECT 2665.730 1051.090 2666.910 1052.270 ;
        RECT 2664.130 1049.490 2665.310 1050.670 ;
        RECT 2665.730 1049.490 2666.910 1050.670 ;
        RECT 2664.130 871.090 2665.310 872.270 ;
        RECT 2665.730 871.090 2666.910 872.270 ;
        RECT 2664.130 869.490 2665.310 870.670 ;
        RECT 2665.730 869.490 2666.910 870.670 ;
        RECT 2664.130 691.090 2665.310 692.270 ;
        RECT 2665.730 691.090 2666.910 692.270 ;
        RECT 2664.130 689.490 2665.310 690.670 ;
        RECT 2665.730 689.490 2666.910 690.670 ;
        RECT 2664.130 511.090 2665.310 512.270 ;
        RECT 2665.730 511.090 2666.910 512.270 ;
        RECT 2664.130 509.490 2665.310 510.670 ;
        RECT 2665.730 509.490 2666.910 510.670 ;
        RECT 2664.130 331.090 2665.310 332.270 ;
        RECT 2665.730 331.090 2666.910 332.270 ;
        RECT 2664.130 329.490 2665.310 330.670 ;
        RECT 2665.730 329.490 2666.910 330.670 ;
        RECT 2664.130 151.090 2665.310 152.270 ;
        RECT 2665.730 151.090 2666.910 152.270 ;
        RECT 2664.130 149.490 2665.310 150.670 ;
        RECT 2665.730 149.490 2666.910 150.670 ;
        RECT 2664.130 -31.710 2665.310 -30.530 ;
        RECT 2665.730 -31.710 2666.910 -30.530 ;
        RECT 2664.130 -33.310 2665.310 -32.130 ;
        RECT 2665.730 -33.310 2666.910 -32.130 ;
        RECT 2844.130 3551.810 2845.310 3552.990 ;
        RECT 2845.730 3551.810 2846.910 3552.990 ;
        RECT 2844.130 3550.210 2845.310 3551.390 ;
        RECT 2845.730 3550.210 2846.910 3551.390 ;
        RECT 2844.130 3391.090 2845.310 3392.270 ;
        RECT 2845.730 3391.090 2846.910 3392.270 ;
        RECT 2844.130 3389.490 2845.310 3390.670 ;
        RECT 2845.730 3389.490 2846.910 3390.670 ;
        RECT 2844.130 3211.090 2845.310 3212.270 ;
        RECT 2845.730 3211.090 2846.910 3212.270 ;
        RECT 2844.130 3209.490 2845.310 3210.670 ;
        RECT 2845.730 3209.490 2846.910 3210.670 ;
        RECT 2844.130 3031.090 2845.310 3032.270 ;
        RECT 2845.730 3031.090 2846.910 3032.270 ;
        RECT 2844.130 3029.490 2845.310 3030.670 ;
        RECT 2845.730 3029.490 2846.910 3030.670 ;
        RECT 2844.130 2851.090 2845.310 2852.270 ;
        RECT 2845.730 2851.090 2846.910 2852.270 ;
        RECT 2844.130 2849.490 2845.310 2850.670 ;
        RECT 2845.730 2849.490 2846.910 2850.670 ;
        RECT 2844.130 2671.090 2845.310 2672.270 ;
        RECT 2845.730 2671.090 2846.910 2672.270 ;
        RECT 2844.130 2669.490 2845.310 2670.670 ;
        RECT 2845.730 2669.490 2846.910 2670.670 ;
        RECT 2844.130 2491.090 2845.310 2492.270 ;
        RECT 2845.730 2491.090 2846.910 2492.270 ;
        RECT 2844.130 2489.490 2845.310 2490.670 ;
        RECT 2845.730 2489.490 2846.910 2490.670 ;
        RECT 2844.130 2311.090 2845.310 2312.270 ;
        RECT 2845.730 2311.090 2846.910 2312.270 ;
        RECT 2844.130 2309.490 2845.310 2310.670 ;
        RECT 2845.730 2309.490 2846.910 2310.670 ;
        RECT 2844.130 2131.090 2845.310 2132.270 ;
        RECT 2845.730 2131.090 2846.910 2132.270 ;
        RECT 2844.130 2129.490 2845.310 2130.670 ;
        RECT 2845.730 2129.490 2846.910 2130.670 ;
        RECT 2844.130 1951.090 2845.310 1952.270 ;
        RECT 2845.730 1951.090 2846.910 1952.270 ;
        RECT 2844.130 1949.490 2845.310 1950.670 ;
        RECT 2845.730 1949.490 2846.910 1950.670 ;
        RECT 2844.130 1771.090 2845.310 1772.270 ;
        RECT 2845.730 1771.090 2846.910 1772.270 ;
        RECT 2844.130 1769.490 2845.310 1770.670 ;
        RECT 2845.730 1769.490 2846.910 1770.670 ;
        RECT 2844.130 1591.090 2845.310 1592.270 ;
        RECT 2845.730 1591.090 2846.910 1592.270 ;
        RECT 2844.130 1589.490 2845.310 1590.670 ;
        RECT 2845.730 1589.490 2846.910 1590.670 ;
        RECT 2844.130 1411.090 2845.310 1412.270 ;
        RECT 2845.730 1411.090 2846.910 1412.270 ;
        RECT 2844.130 1409.490 2845.310 1410.670 ;
        RECT 2845.730 1409.490 2846.910 1410.670 ;
        RECT 2844.130 1231.090 2845.310 1232.270 ;
        RECT 2845.730 1231.090 2846.910 1232.270 ;
        RECT 2844.130 1229.490 2845.310 1230.670 ;
        RECT 2845.730 1229.490 2846.910 1230.670 ;
        RECT 2844.130 1051.090 2845.310 1052.270 ;
        RECT 2845.730 1051.090 2846.910 1052.270 ;
        RECT 2844.130 1049.490 2845.310 1050.670 ;
        RECT 2845.730 1049.490 2846.910 1050.670 ;
        RECT 2844.130 871.090 2845.310 872.270 ;
        RECT 2845.730 871.090 2846.910 872.270 ;
        RECT 2844.130 869.490 2845.310 870.670 ;
        RECT 2845.730 869.490 2846.910 870.670 ;
        RECT 2844.130 691.090 2845.310 692.270 ;
        RECT 2845.730 691.090 2846.910 692.270 ;
        RECT 2844.130 689.490 2845.310 690.670 ;
        RECT 2845.730 689.490 2846.910 690.670 ;
        RECT 2844.130 511.090 2845.310 512.270 ;
        RECT 2845.730 511.090 2846.910 512.270 ;
        RECT 2844.130 509.490 2845.310 510.670 ;
        RECT 2845.730 509.490 2846.910 510.670 ;
        RECT 2844.130 331.090 2845.310 332.270 ;
        RECT 2845.730 331.090 2846.910 332.270 ;
        RECT 2844.130 329.490 2845.310 330.670 ;
        RECT 2845.730 329.490 2846.910 330.670 ;
        RECT 2844.130 151.090 2845.310 152.270 ;
        RECT 2845.730 151.090 2846.910 152.270 ;
        RECT 2844.130 149.490 2845.310 150.670 ;
        RECT 2845.730 149.490 2846.910 150.670 ;
        RECT 2844.130 -31.710 2845.310 -30.530 ;
        RECT 2845.730 -31.710 2846.910 -30.530 ;
        RECT 2844.130 -33.310 2845.310 -32.130 ;
        RECT 2845.730 -33.310 2846.910 -32.130 ;
        RECT 2955.510 3551.810 2956.690 3552.990 ;
        RECT 2957.110 3551.810 2958.290 3552.990 ;
        RECT 2955.510 3550.210 2956.690 3551.390 ;
        RECT 2957.110 3550.210 2958.290 3551.390 ;
        RECT 2955.510 3391.090 2956.690 3392.270 ;
        RECT 2957.110 3391.090 2958.290 3392.270 ;
        RECT 2955.510 3389.490 2956.690 3390.670 ;
        RECT 2957.110 3389.490 2958.290 3390.670 ;
        RECT 2955.510 3211.090 2956.690 3212.270 ;
        RECT 2957.110 3211.090 2958.290 3212.270 ;
        RECT 2955.510 3209.490 2956.690 3210.670 ;
        RECT 2957.110 3209.490 2958.290 3210.670 ;
        RECT 2955.510 3031.090 2956.690 3032.270 ;
        RECT 2957.110 3031.090 2958.290 3032.270 ;
        RECT 2955.510 3029.490 2956.690 3030.670 ;
        RECT 2957.110 3029.490 2958.290 3030.670 ;
        RECT 2955.510 2851.090 2956.690 2852.270 ;
        RECT 2957.110 2851.090 2958.290 2852.270 ;
        RECT 2955.510 2849.490 2956.690 2850.670 ;
        RECT 2957.110 2849.490 2958.290 2850.670 ;
        RECT 2955.510 2671.090 2956.690 2672.270 ;
        RECT 2957.110 2671.090 2958.290 2672.270 ;
        RECT 2955.510 2669.490 2956.690 2670.670 ;
        RECT 2957.110 2669.490 2958.290 2670.670 ;
        RECT 2955.510 2491.090 2956.690 2492.270 ;
        RECT 2957.110 2491.090 2958.290 2492.270 ;
        RECT 2955.510 2489.490 2956.690 2490.670 ;
        RECT 2957.110 2489.490 2958.290 2490.670 ;
        RECT 2955.510 2311.090 2956.690 2312.270 ;
        RECT 2957.110 2311.090 2958.290 2312.270 ;
        RECT 2955.510 2309.490 2956.690 2310.670 ;
        RECT 2957.110 2309.490 2958.290 2310.670 ;
        RECT 2955.510 2131.090 2956.690 2132.270 ;
        RECT 2957.110 2131.090 2958.290 2132.270 ;
        RECT 2955.510 2129.490 2956.690 2130.670 ;
        RECT 2957.110 2129.490 2958.290 2130.670 ;
        RECT 2955.510 1951.090 2956.690 1952.270 ;
        RECT 2957.110 1951.090 2958.290 1952.270 ;
        RECT 2955.510 1949.490 2956.690 1950.670 ;
        RECT 2957.110 1949.490 2958.290 1950.670 ;
        RECT 2955.510 1771.090 2956.690 1772.270 ;
        RECT 2957.110 1771.090 2958.290 1772.270 ;
        RECT 2955.510 1769.490 2956.690 1770.670 ;
        RECT 2957.110 1769.490 2958.290 1770.670 ;
        RECT 2955.510 1591.090 2956.690 1592.270 ;
        RECT 2957.110 1591.090 2958.290 1592.270 ;
        RECT 2955.510 1589.490 2956.690 1590.670 ;
        RECT 2957.110 1589.490 2958.290 1590.670 ;
        RECT 2955.510 1411.090 2956.690 1412.270 ;
        RECT 2957.110 1411.090 2958.290 1412.270 ;
        RECT 2955.510 1409.490 2956.690 1410.670 ;
        RECT 2957.110 1409.490 2958.290 1410.670 ;
        RECT 2955.510 1231.090 2956.690 1232.270 ;
        RECT 2957.110 1231.090 2958.290 1232.270 ;
        RECT 2955.510 1229.490 2956.690 1230.670 ;
        RECT 2957.110 1229.490 2958.290 1230.670 ;
        RECT 2955.510 1051.090 2956.690 1052.270 ;
        RECT 2957.110 1051.090 2958.290 1052.270 ;
        RECT 2955.510 1049.490 2956.690 1050.670 ;
        RECT 2957.110 1049.490 2958.290 1050.670 ;
        RECT 2955.510 871.090 2956.690 872.270 ;
        RECT 2957.110 871.090 2958.290 872.270 ;
        RECT 2955.510 869.490 2956.690 870.670 ;
        RECT 2957.110 869.490 2958.290 870.670 ;
        RECT 2955.510 691.090 2956.690 692.270 ;
        RECT 2957.110 691.090 2958.290 692.270 ;
        RECT 2955.510 689.490 2956.690 690.670 ;
        RECT 2957.110 689.490 2958.290 690.670 ;
        RECT 2955.510 511.090 2956.690 512.270 ;
        RECT 2957.110 511.090 2958.290 512.270 ;
        RECT 2955.510 509.490 2956.690 510.670 ;
        RECT 2957.110 509.490 2958.290 510.670 ;
        RECT 2955.510 331.090 2956.690 332.270 ;
        RECT 2957.110 331.090 2958.290 332.270 ;
        RECT 2955.510 329.490 2956.690 330.670 ;
        RECT 2957.110 329.490 2958.290 330.670 ;
        RECT 2955.510 151.090 2956.690 152.270 ;
        RECT 2957.110 151.090 2958.290 152.270 ;
        RECT 2955.510 149.490 2956.690 150.670 ;
        RECT 2957.110 149.490 2958.290 150.670 ;
        RECT 2955.510 -31.710 2956.690 -30.530 ;
        RECT 2957.110 -31.710 2958.290 -30.530 ;
        RECT 2955.510 -33.310 2956.690 -32.130 ;
        RECT 2957.110 -33.310 2958.290 -32.130 ;
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
        RECT -43.630 3389.330 2963.250 3392.430 ;
        RECT -43.630 3209.330 2963.250 3212.430 ;
        RECT -43.630 3029.330 2963.250 3032.430 ;
        RECT -43.630 2849.330 2963.250 2852.430 ;
        RECT -43.630 2669.330 2963.250 2672.430 ;
        RECT -43.630 2489.330 2963.250 2492.430 ;
        RECT -43.630 2309.330 2963.250 2312.430 ;
        RECT -43.630 2129.330 2963.250 2132.430 ;
        RECT -43.630 1949.330 2963.250 1952.430 ;
        RECT -43.630 1769.330 2963.250 1772.430 ;
        RECT -43.630 1589.330 2963.250 1592.430 ;
        RECT -43.630 1409.330 2963.250 1412.430 ;
        RECT -43.630 1229.330 2963.250 1232.430 ;
        RECT -43.630 1049.330 2963.250 1052.430 ;
        RECT -43.630 869.330 2963.250 872.430 ;
        RECT -43.630 689.330 2963.250 692.430 ;
        RECT -43.630 509.330 2963.250 512.430 ;
        RECT -43.630 329.330 2963.250 332.430 ;
        RECT -43.630 149.330 2963.250 152.430 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
        RECT 121.470 -38.270 124.570 3557.950 ;
        RECT 301.470 -38.270 304.570 3557.950 ;
        RECT 481.470 810.000 484.570 3557.950 ;
        RECT 661.470 810.000 664.570 3557.950 ;
        RECT 481.470 -38.270 484.570 490.000 ;
        RECT 661.470 -38.270 664.570 490.000 ;
        RECT 841.470 -38.270 844.570 3557.950 ;
        RECT 1021.470 -38.270 1024.570 3557.950 ;
        RECT 1201.470 -38.270 1204.570 3557.950 ;
        RECT 1381.470 -38.270 1384.570 3557.950 ;
        RECT 1561.470 -38.270 1564.570 3557.950 ;
        RECT 1741.470 -38.270 1744.570 3557.950 ;
        RECT 1921.470 -38.270 1924.570 3557.950 ;
        RECT 2101.470 -38.270 2104.570 3557.950 ;
        RECT 2281.470 -38.270 2284.570 3557.950 ;
        RECT 2461.470 -38.270 2464.570 3557.950 ;
        RECT 2641.470 -38.270 2644.570 3557.950 ;
        RECT 2821.470 -38.270 2824.570 3557.950 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
      LAYER via4 ;
        RECT -33.870 3547.010 -32.690 3548.190 ;
        RECT -32.270 3547.010 -31.090 3548.190 ;
        RECT -33.870 3545.410 -32.690 3546.590 ;
        RECT -32.270 3545.410 -31.090 3546.590 ;
        RECT -33.870 3368.590 -32.690 3369.770 ;
        RECT -32.270 3368.590 -31.090 3369.770 ;
        RECT -33.870 3366.990 -32.690 3368.170 ;
        RECT -32.270 3366.990 -31.090 3368.170 ;
        RECT -33.870 3188.590 -32.690 3189.770 ;
        RECT -32.270 3188.590 -31.090 3189.770 ;
        RECT -33.870 3186.990 -32.690 3188.170 ;
        RECT -32.270 3186.990 -31.090 3188.170 ;
        RECT -33.870 3008.590 -32.690 3009.770 ;
        RECT -32.270 3008.590 -31.090 3009.770 ;
        RECT -33.870 3006.990 -32.690 3008.170 ;
        RECT -32.270 3006.990 -31.090 3008.170 ;
        RECT -33.870 2828.590 -32.690 2829.770 ;
        RECT -32.270 2828.590 -31.090 2829.770 ;
        RECT -33.870 2826.990 -32.690 2828.170 ;
        RECT -32.270 2826.990 -31.090 2828.170 ;
        RECT -33.870 2648.590 -32.690 2649.770 ;
        RECT -32.270 2648.590 -31.090 2649.770 ;
        RECT -33.870 2646.990 -32.690 2648.170 ;
        RECT -32.270 2646.990 -31.090 2648.170 ;
        RECT -33.870 2468.590 -32.690 2469.770 ;
        RECT -32.270 2468.590 -31.090 2469.770 ;
        RECT -33.870 2466.990 -32.690 2468.170 ;
        RECT -32.270 2466.990 -31.090 2468.170 ;
        RECT -33.870 2288.590 -32.690 2289.770 ;
        RECT -32.270 2288.590 -31.090 2289.770 ;
        RECT -33.870 2286.990 -32.690 2288.170 ;
        RECT -32.270 2286.990 -31.090 2288.170 ;
        RECT -33.870 2108.590 -32.690 2109.770 ;
        RECT -32.270 2108.590 -31.090 2109.770 ;
        RECT -33.870 2106.990 -32.690 2108.170 ;
        RECT -32.270 2106.990 -31.090 2108.170 ;
        RECT -33.870 1928.590 -32.690 1929.770 ;
        RECT -32.270 1928.590 -31.090 1929.770 ;
        RECT -33.870 1926.990 -32.690 1928.170 ;
        RECT -32.270 1926.990 -31.090 1928.170 ;
        RECT -33.870 1748.590 -32.690 1749.770 ;
        RECT -32.270 1748.590 -31.090 1749.770 ;
        RECT -33.870 1746.990 -32.690 1748.170 ;
        RECT -32.270 1746.990 -31.090 1748.170 ;
        RECT -33.870 1568.590 -32.690 1569.770 ;
        RECT -32.270 1568.590 -31.090 1569.770 ;
        RECT -33.870 1566.990 -32.690 1568.170 ;
        RECT -32.270 1566.990 -31.090 1568.170 ;
        RECT -33.870 1388.590 -32.690 1389.770 ;
        RECT -32.270 1388.590 -31.090 1389.770 ;
        RECT -33.870 1386.990 -32.690 1388.170 ;
        RECT -32.270 1386.990 -31.090 1388.170 ;
        RECT -33.870 1208.590 -32.690 1209.770 ;
        RECT -32.270 1208.590 -31.090 1209.770 ;
        RECT -33.870 1206.990 -32.690 1208.170 ;
        RECT -32.270 1206.990 -31.090 1208.170 ;
        RECT -33.870 1028.590 -32.690 1029.770 ;
        RECT -32.270 1028.590 -31.090 1029.770 ;
        RECT -33.870 1026.990 -32.690 1028.170 ;
        RECT -32.270 1026.990 -31.090 1028.170 ;
        RECT -33.870 848.590 -32.690 849.770 ;
        RECT -32.270 848.590 -31.090 849.770 ;
        RECT -33.870 846.990 -32.690 848.170 ;
        RECT -32.270 846.990 -31.090 848.170 ;
        RECT -33.870 668.590 -32.690 669.770 ;
        RECT -32.270 668.590 -31.090 669.770 ;
        RECT -33.870 666.990 -32.690 668.170 ;
        RECT -32.270 666.990 -31.090 668.170 ;
        RECT -33.870 488.590 -32.690 489.770 ;
        RECT -32.270 488.590 -31.090 489.770 ;
        RECT -33.870 486.990 -32.690 488.170 ;
        RECT -32.270 486.990 -31.090 488.170 ;
        RECT -33.870 308.590 -32.690 309.770 ;
        RECT -32.270 308.590 -31.090 309.770 ;
        RECT -33.870 306.990 -32.690 308.170 ;
        RECT -32.270 306.990 -31.090 308.170 ;
        RECT -33.870 128.590 -32.690 129.770 ;
        RECT -32.270 128.590 -31.090 129.770 ;
        RECT -33.870 126.990 -32.690 128.170 ;
        RECT -32.270 126.990 -31.090 128.170 ;
        RECT -33.870 -26.910 -32.690 -25.730 ;
        RECT -32.270 -26.910 -31.090 -25.730 ;
        RECT -33.870 -28.510 -32.690 -27.330 ;
        RECT -32.270 -28.510 -31.090 -27.330 ;
        RECT 121.630 3547.010 122.810 3548.190 ;
        RECT 123.230 3547.010 124.410 3548.190 ;
        RECT 121.630 3545.410 122.810 3546.590 ;
        RECT 123.230 3545.410 124.410 3546.590 ;
        RECT 121.630 3368.590 122.810 3369.770 ;
        RECT 123.230 3368.590 124.410 3369.770 ;
        RECT 121.630 3366.990 122.810 3368.170 ;
        RECT 123.230 3366.990 124.410 3368.170 ;
        RECT 121.630 3188.590 122.810 3189.770 ;
        RECT 123.230 3188.590 124.410 3189.770 ;
        RECT 121.630 3186.990 122.810 3188.170 ;
        RECT 123.230 3186.990 124.410 3188.170 ;
        RECT 121.630 3008.590 122.810 3009.770 ;
        RECT 123.230 3008.590 124.410 3009.770 ;
        RECT 121.630 3006.990 122.810 3008.170 ;
        RECT 123.230 3006.990 124.410 3008.170 ;
        RECT 121.630 2828.590 122.810 2829.770 ;
        RECT 123.230 2828.590 124.410 2829.770 ;
        RECT 121.630 2826.990 122.810 2828.170 ;
        RECT 123.230 2826.990 124.410 2828.170 ;
        RECT 121.630 2648.590 122.810 2649.770 ;
        RECT 123.230 2648.590 124.410 2649.770 ;
        RECT 121.630 2646.990 122.810 2648.170 ;
        RECT 123.230 2646.990 124.410 2648.170 ;
        RECT 121.630 2468.590 122.810 2469.770 ;
        RECT 123.230 2468.590 124.410 2469.770 ;
        RECT 121.630 2466.990 122.810 2468.170 ;
        RECT 123.230 2466.990 124.410 2468.170 ;
        RECT 121.630 2288.590 122.810 2289.770 ;
        RECT 123.230 2288.590 124.410 2289.770 ;
        RECT 121.630 2286.990 122.810 2288.170 ;
        RECT 123.230 2286.990 124.410 2288.170 ;
        RECT 121.630 2108.590 122.810 2109.770 ;
        RECT 123.230 2108.590 124.410 2109.770 ;
        RECT 121.630 2106.990 122.810 2108.170 ;
        RECT 123.230 2106.990 124.410 2108.170 ;
        RECT 121.630 1928.590 122.810 1929.770 ;
        RECT 123.230 1928.590 124.410 1929.770 ;
        RECT 121.630 1926.990 122.810 1928.170 ;
        RECT 123.230 1926.990 124.410 1928.170 ;
        RECT 121.630 1748.590 122.810 1749.770 ;
        RECT 123.230 1748.590 124.410 1749.770 ;
        RECT 121.630 1746.990 122.810 1748.170 ;
        RECT 123.230 1746.990 124.410 1748.170 ;
        RECT 121.630 1568.590 122.810 1569.770 ;
        RECT 123.230 1568.590 124.410 1569.770 ;
        RECT 121.630 1566.990 122.810 1568.170 ;
        RECT 123.230 1566.990 124.410 1568.170 ;
        RECT 121.630 1388.590 122.810 1389.770 ;
        RECT 123.230 1388.590 124.410 1389.770 ;
        RECT 121.630 1386.990 122.810 1388.170 ;
        RECT 123.230 1386.990 124.410 1388.170 ;
        RECT 121.630 1208.590 122.810 1209.770 ;
        RECT 123.230 1208.590 124.410 1209.770 ;
        RECT 121.630 1206.990 122.810 1208.170 ;
        RECT 123.230 1206.990 124.410 1208.170 ;
        RECT 121.630 1028.590 122.810 1029.770 ;
        RECT 123.230 1028.590 124.410 1029.770 ;
        RECT 121.630 1026.990 122.810 1028.170 ;
        RECT 123.230 1026.990 124.410 1028.170 ;
        RECT 121.630 848.590 122.810 849.770 ;
        RECT 123.230 848.590 124.410 849.770 ;
        RECT 121.630 846.990 122.810 848.170 ;
        RECT 123.230 846.990 124.410 848.170 ;
        RECT 121.630 668.590 122.810 669.770 ;
        RECT 123.230 668.590 124.410 669.770 ;
        RECT 121.630 666.990 122.810 668.170 ;
        RECT 123.230 666.990 124.410 668.170 ;
        RECT 121.630 488.590 122.810 489.770 ;
        RECT 123.230 488.590 124.410 489.770 ;
        RECT 121.630 486.990 122.810 488.170 ;
        RECT 123.230 486.990 124.410 488.170 ;
        RECT 121.630 308.590 122.810 309.770 ;
        RECT 123.230 308.590 124.410 309.770 ;
        RECT 121.630 306.990 122.810 308.170 ;
        RECT 123.230 306.990 124.410 308.170 ;
        RECT 121.630 128.590 122.810 129.770 ;
        RECT 123.230 128.590 124.410 129.770 ;
        RECT 121.630 126.990 122.810 128.170 ;
        RECT 123.230 126.990 124.410 128.170 ;
        RECT 121.630 -26.910 122.810 -25.730 ;
        RECT 123.230 -26.910 124.410 -25.730 ;
        RECT 121.630 -28.510 122.810 -27.330 ;
        RECT 123.230 -28.510 124.410 -27.330 ;
        RECT 301.630 3547.010 302.810 3548.190 ;
        RECT 303.230 3547.010 304.410 3548.190 ;
        RECT 301.630 3545.410 302.810 3546.590 ;
        RECT 303.230 3545.410 304.410 3546.590 ;
        RECT 301.630 3368.590 302.810 3369.770 ;
        RECT 303.230 3368.590 304.410 3369.770 ;
        RECT 301.630 3366.990 302.810 3368.170 ;
        RECT 303.230 3366.990 304.410 3368.170 ;
        RECT 301.630 3188.590 302.810 3189.770 ;
        RECT 303.230 3188.590 304.410 3189.770 ;
        RECT 301.630 3186.990 302.810 3188.170 ;
        RECT 303.230 3186.990 304.410 3188.170 ;
        RECT 301.630 3008.590 302.810 3009.770 ;
        RECT 303.230 3008.590 304.410 3009.770 ;
        RECT 301.630 3006.990 302.810 3008.170 ;
        RECT 303.230 3006.990 304.410 3008.170 ;
        RECT 301.630 2828.590 302.810 2829.770 ;
        RECT 303.230 2828.590 304.410 2829.770 ;
        RECT 301.630 2826.990 302.810 2828.170 ;
        RECT 303.230 2826.990 304.410 2828.170 ;
        RECT 301.630 2648.590 302.810 2649.770 ;
        RECT 303.230 2648.590 304.410 2649.770 ;
        RECT 301.630 2646.990 302.810 2648.170 ;
        RECT 303.230 2646.990 304.410 2648.170 ;
        RECT 301.630 2468.590 302.810 2469.770 ;
        RECT 303.230 2468.590 304.410 2469.770 ;
        RECT 301.630 2466.990 302.810 2468.170 ;
        RECT 303.230 2466.990 304.410 2468.170 ;
        RECT 301.630 2288.590 302.810 2289.770 ;
        RECT 303.230 2288.590 304.410 2289.770 ;
        RECT 301.630 2286.990 302.810 2288.170 ;
        RECT 303.230 2286.990 304.410 2288.170 ;
        RECT 301.630 2108.590 302.810 2109.770 ;
        RECT 303.230 2108.590 304.410 2109.770 ;
        RECT 301.630 2106.990 302.810 2108.170 ;
        RECT 303.230 2106.990 304.410 2108.170 ;
        RECT 301.630 1928.590 302.810 1929.770 ;
        RECT 303.230 1928.590 304.410 1929.770 ;
        RECT 301.630 1926.990 302.810 1928.170 ;
        RECT 303.230 1926.990 304.410 1928.170 ;
        RECT 301.630 1748.590 302.810 1749.770 ;
        RECT 303.230 1748.590 304.410 1749.770 ;
        RECT 301.630 1746.990 302.810 1748.170 ;
        RECT 303.230 1746.990 304.410 1748.170 ;
        RECT 301.630 1568.590 302.810 1569.770 ;
        RECT 303.230 1568.590 304.410 1569.770 ;
        RECT 301.630 1566.990 302.810 1568.170 ;
        RECT 303.230 1566.990 304.410 1568.170 ;
        RECT 301.630 1388.590 302.810 1389.770 ;
        RECT 303.230 1388.590 304.410 1389.770 ;
        RECT 301.630 1386.990 302.810 1388.170 ;
        RECT 303.230 1386.990 304.410 1388.170 ;
        RECT 301.630 1208.590 302.810 1209.770 ;
        RECT 303.230 1208.590 304.410 1209.770 ;
        RECT 301.630 1206.990 302.810 1208.170 ;
        RECT 303.230 1206.990 304.410 1208.170 ;
        RECT 301.630 1028.590 302.810 1029.770 ;
        RECT 303.230 1028.590 304.410 1029.770 ;
        RECT 301.630 1026.990 302.810 1028.170 ;
        RECT 303.230 1026.990 304.410 1028.170 ;
        RECT 301.630 848.590 302.810 849.770 ;
        RECT 303.230 848.590 304.410 849.770 ;
        RECT 301.630 846.990 302.810 848.170 ;
        RECT 303.230 846.990 304.410 848.170 ;
        RECT 481.630 3547.010 482.810 3548.190 ;
        RECT 483.230 3547.010 484.410 3548.190 ;
        RECT 481.630 3545.410 482.810 3546.590 ;
        RECT 483.230 3545.410 484.410 3546.590 ;
        RECT 481.630 3368.590 482.810 3369.770 ;
        RECT 483.230 3368.590 484.410 3369.770 ;
        RECT 481.630 3366.990 482.810 3368.170 ;
        RECT 483.230 3366.990 484.410 3368.170 ;
        RECT 481.630 3188.590 482.810 3189.770 ;
        RECT 483.230 3188.590 484.410 3189.770 ;
        RECT 481.630 3186.990 482.810 3188.170 ;
        RECT 483.230 3186.990 484.410 3188.170 ;
        RECT 481.630 3008.590 482.810 3009.770 ;
        RECT 483.230 3008.590 484.410 3009.770 ;
        RECT 481.630 3006.990 482.810 3008.170 ;
        RECT 483.230 3006.990 484.410 3008.170 ;
        RECT 481.630 2828.590 482.810 2829.770 ;
        RECT 483.230 2828.590 484.410 2829.770 ;
        RECT 481.630 2826.990 482.810 2828.170 ;
        RECT 483.230 2826.990 484.410 2828.170 ;
        RECT 481.630 2648.590 482.810 2649.770 ;
        RECT 483.230 2648.590 484.410 2649.770 ;
        RECT 481.630 2646.990 482.810 2648.170 ;
        RECT 483.230 2646.990 484.410 2648.170 ;
        RECT 481.630 2468.590 482.810 2469.770 ;
        RECT 483.230 2468.590 484.410 2469.770 ;
        RECT 481.630 2466.990 482.810 2468.170 ;
        RECT 483.230 2466.990 484.410 2468.170 ;
        RECT 481.630 2288.590 482.810 2289.770 ;
        RECT 483.230 2288.590 484.410 2289.770 ;
        RECT 481.630 2286.990 482.810 2288.170 ;
        RECT 483.230 2286.990 484.410 2288.170 ;
        RECT 481.630 2108.590 482.810 2109.770 ;
        RECT 483.230 2108.590 484.410 2109.770 ;
        RECT 481.630 2106.990 482.810 2108.170 ;
        RECT 483.230 2106.990 484.410 2108.170 ;
        RECT 481.630 1928.590 482.810 1929.770 ;
        RECT 483.230 1928.590 484.410 1929.770 ;
        RECT 481.630 1926.990 482.810 1928.170 ;
        RECT 483.230 1926.990 484.410 1928.170 ;
        RECT 481.630 1748.590 482.810 1749.770 ;
        RECT 483.230 1748.590 484.410 1749.770 ;
        RECT 481.630 1746.990 482.810 1748.170 ;
        RECT 483.230 1746.990 484.410 1748.170 ;
        RECT 481.630 1568.590 482.810 1569.770 ;
        RECT 483.230 1568.590 484.410 1569.770 ;
        RECT 481.630 1566.990 482.810 1568.170 ;
        RECT 483.230 1566.990 484.410 1568.170 ;
        RECT 481.630 1388.590 482.810 1389.770 ;
        RECT 483.230 1388.590 484.410 1389.770 ;
        RECT 481.630 1386.990 482.810 1388.170 ;
        RECT 483.230 1386.990 484.410 1388.170 ;
        RECT 481.630 1208.590 482.810 1209.770 ;
        RECT 483.230 1208.590 484.410 1209.770 ;
        RECT 481.630 1206.990 482.810 1208.170 ;
        RECT 483.230 1206.990 484.410 1208.170 ;
        RECT 481.630 1028.590 482.810 1029.770 ;
        RECT 483.230 1028.590 484.410 1029.770 ;
        RECT 481.630 1026.990 482.810 1028.170 ;
        RECT 483.230 1026.990 484.410 1028.170 ;
        RECT 481.630 848.590 482.810 849.770 ;
        RECT 483.230 848.590 484.410 849.770 ;
        RECT 481.630 846.990 482.810 848.170 ;
        RECT 483.230 846.990 484.410 848.170 ;
        RECT 661.630 3547.010 662.810 3548.190 ;
        RECT 663.230 3547.010 664.410 3548.190 ;
        RECT 661.630 3545.410 662.810 3546.590 ;
        RECT 663.230 3545.410 664.410 3546.590 ;
        RECT 661.630 3368.590 662.810 3369.770 ;
        RECT 663.230 3368.590 664.410 3369.770 ;
        RECT 661.630 3366.990 662.810 3368.170 ;
        RECT 663.230 3366.990 664.410 3368.170 ;
        RECT 661.630 3188.590 662.810 3189.770 ;
        RECT 663.230 3188.590 664.410 3189.770 ;
        RECT 661.630 3186.990 662.810 3188.170 ;
        RECT 663.230 3186.990 664.410 3188.170 ;
        RECT 661.630 3008.590 662.810 3009.770 ;
        RECT 663.230 3008.590 664.410 3009.770 ;
        RECT 661.630 3006.990 662.810 3008.170 ;
        RECT 663.230 3006.990 664.410 3008.170 ;
        RECT 661.630 2828.590 662.810 2829.770 ;
        RECT 663.230 2828.590 664.410 2829.770 ;
        RECT 661.630 2826.990 662.810 2828.170 ;
        RECT 663.230 2826.990 664.410 2828.170 ;
        RECT 661.630 2648.590 662.810 2649.770 ;
        RECT 663.230 2648.590 664.410 2649.770 ;
        RECT 661.630 2646.990 662.810 2648.170 ;
        RECT 663.230 2646.990 664.410 2648.170 ;
        RECT 661.630 2468.590 662.810 2469.770 ;
        RECT 663.230 2468.590 664.410 2469.770 ;
        RECT 661.630 2466.990 662.810 2468.170 ;
        RECT 663.230 2466.990 664.410 2468.170 ;
        RECT 661.630 2288.590 662.810 2289.770 ;
        RECT 663.230 2288.590 664.410 2289.770 ;
        RECT 661.630 2286.990 662.810 2288.170 ;
        RECT 663.230 2286.990 664.410 2288.170 ;
        RECT 661.630 2108.590 662.810 2109.770 ;
        RECT 663.230 2108.590 664.410 2109.770 ;
        RECT 661.630 2106.990 662.810 2108.170 ;
        RECT 663.230 2106.990 664.410 2108.170 ;
        RECT 661.630 1928.590 662.810 1929.770 ;
        RECT 663.230 1928.590 664.410 1929.770 ;
        RECT 661.630 1926.990 662.810 1928.170 ;
        RECT 663.230 1926.990 664.410 1928.170 ;
        RECT 661.630 1748.590 662.810 1749.770 ;
        RECT 663.230 1748.590 664.410 1749.770 ;
        RECT 661.630 1746.990 662.810 1748.170 ;
        RECT 663.230 1746.990 664.410 1748.170 ;
        RECT 661.630 1568.590 662.810 1569.770 ;
        RECT 663.230 1568.590 664.410 1569.770 ;
        RECT 661.630 1566.990 662.810 1568.170 ;
        RECT 663.230 1566.990 664.410 1568.170 ;
        RECT 661.630 1388.590 662.810 1389.770 ;
        RECT 663.230 1388.590 664.410 1389.770 ;
        RECT 661.630 1386.990 662.810 1388.170 ;
        RECT 663.230 1386.990 664.410 1388.170 ;
        RECT 661.630 1208.590 662.810 1209.770 ;
        RECT 663.230 1208.590 664.410 1209.770 ;
        RECT 661.630 1206.990 662.810 1208.170 ;
        RECT 663.230 1206.990 664.410 1208.170 ;
        RECT 661.630 1028.590 662.810 1029.770 ;
        RECT 663.230 1028.590 664.410 1029.770 ;
        RECT 661.630 1026.990 662.810 1028.170 ;
        RECT 663.230 1026.990 664.410 1028.170 ;
        RECT 661.630 848.590 662.810 849.770 ;
        RECT 663.230 848.590 664.410 849.770 ;
        RECT 661.630 846.990 662.810 848.170 ;
        RECT 663.230 846.990 664.410 848.170 ;
        RECT 841.630 3547.010 842.810 3548.190 ;
        RECT 843.230 3547.010 844.410 3548.190 ;
        RECT 841.630 3545.410 842.810 3546.590 ;
        RECT 843.230 3545.410 844.410 3546.590 ;
        RECT 841.630 3368.590 842.810 3369.770 ;
        RECT 843.230 3368.590 844.410 3369.770 ;
        RECT 841.630 3366.990 842.810 3368.170 ;
        RECT 843.230 3366.990 844.410 3368.170 ;
        RECT 841.630 3188.590 842.810 3189.770 ;
        RECT 843.230 3188.590 844.410 3189.770 ;
        RECT 841.630 3186.990 842.810 3188.170 ;
        RECT 843.230 3186.990 844.410 3188.170 ;
        RECT 841.630 3008.590 842.810 3009.770 ;
        RECT 843.230 3008.590 844.410 3009.770 ;
        RECT 841.630 3006.990 842.810 3008.170 ;
        RECT 843.230 3006.990 844.410 3008.170 ;
        RECT 841.630 2828.590 842.810 2829.770 ;
        RECT 843.230 2828.590 844.410 2829.770 ;
        RECT 841.630 2826.990 842.810 2828.170 ;
        RECT 843.230 2826.990 844.410 2828.170 ;
        RECT 841.630 2648.590 842.810 2649.770 ;
        RECT 843.230 2648.590 844.410 2649.770 ;
        RECT 841.630 2646.990 842.810 2648.170 ;
        RECT 843.230 2646.990 844.410 2648.170 ;
        RECT 841.630 2468.590 842.810 2469.770 ;
        RECT 843.230 2468.590 844.410 2469.770 ;
        RECT 841.630 2466.990 842.810 2468.170 ;
        RECT 843.230 2466.990 844.410 2468.170 ;
        RECT 841.630 2288.590 842.810 2289.770 ;
        RECT 843.230 2288.590 844.410 2289.770 ;
        RECT 841.630 2286.990 842.810 2288.170 ;
        RECT 843.230 2286.990 844.410 2288.170 ;
        RECT 841.630 2108.590 842.810 2109.770 ;
        RECT 843.230 2108.590 844.410 2109.770 ;
        RECT 841.630 2106.990 842.810 2108.170 ;
        RECT 843.230 2106.990 844.410 2108.170 ;
        RECT 841.630 1928.590 842.810 1929.770 ;
        RECT 843.230 1928.590 844.410 1929.770 ;
        RECT 841.630 1926.990 842.810 1928.170 ;
        RECT 843.230 1926.990 844.410 1928.170 ;
        RECT 841.630 1748.590 842.810 1749.770 ;
        RECT 843.230 1748.590 844.410 1749.770 ;
        RECT 841.630 1746.990 842.810 1748.170 ;
        RECT 843.230 1746.990 844.410 1748.170 ;
        RECT 841.630 1568.590 842.810 1569.770 ;
        RECT 843.230 1568.590 844.410 1569.770 ;
        RECT 841.630 1566.990 842.810 1568.170 ;
        RECT 843.230 1566.990 844.410 1568.170 ;
        RECT 841.630 1388.590 842.810 1389.770 ;
        RECT 843.230 1388.590 844.410 1389.770 ;
        RECT 841.630 1386.990 842.810 1388.170 ;
        RECT 843.230 1386.990 844.410 1388.170 ;
        RECT 841.630 1208.590 842.810 1209.770 ;
        RECT 843.230 1208.590 844.410 1209.770 ;
        RECT 841.630 1206.990 842.810 1208.170 ;
        RECT 843.230 1206.990 844.410 1208.170 ;
        RECT 841.630 1028.590 842.810 1029.770 ;
        RECT 843.230 1028.590 844.410 1029.770 ;
        RECT 841.630 1026.990 842.810 1028.170 ;
        RECT 843.230 1026.990 844.410 1028.170 ;
        RECT 841.630 848.590 842.810 849.770 ;
        RECT 843.230 848.590 844.410 849.770 ;
        RECT 841.630 846.990 842.810 848.170 ;
        RECT 843.230 846.990 844.410 848.170 ;
        RECT 301.630 668.590 302.810 669.770 ;
        RECT 303.230 668.590 304.410 669.770 ;
        RECT 301.630 666.990 302.810 668.170 ;
        RECT 303.230 666.990 304.410 668.170 ;
        RECT 841.630 668.590 842.810 669.770 ;
        RECT 843.230 668.590 844.410 669.770 ;
        RECT 841.630 666.990 842.810 668.170 ;
        RECT 843.230 666.990 844.410 668.170 ;
        RECT 301.630 488.590 302.810 489.770 ;
        RECT 303.230 488.590 304.410 489.770 ;
        RECT 301.630 486.990 302.810 488.170 ;
        RECT 303.230 486.990 304.410 488.170 ;
        RECT 301.630 308.590 302.810 309.770 ;
        RECT 303.230 308.590 304.410 309.770 ;
        RECT 301.630 306.990 302.810 308.170 ;
        RECT 303.230 306.990 304.410 308.170 ;
        RECT 301.630 128.590 302.810 129.770 ;
        RECT 303.230 128.590 304.410 129.770 ;
        RECT 301.630 126.990 302.810 128.170 ;
        RECT 303.230 126.990 304.410 128.170 ;
        RECT 301.630 -26.910 302.810 -25.730 ;
        RECT 303.230 -26.910 304.410 -25.730 ;
        RECT 301.630 -28.510 302.810 -27.330 ;
        RECT 303.230 -28.510 304.410 -27.330 ;
        RECT 481.630 488.590 482.810 489.770 ;
        RECT 483.230 488.590 484.410 489.770 ;
        RECT 481.630 486.990 482.810 488.170 ;
        RECT 483.230 486.990 484.410 488.170 ;
        RECT 481.630 308.590 482.810 309.770 ;
        RECT 483.230 308.590 484.410 309.770 ;
        RECT 481.630 306.990 482.810 308.170 ;
        RECT 483.230 306.990 484.410 308.170 ;
        RECT 481.630 128.590 482.810 129.770 ;
        RECT 483.230 128.590 484.410 129.770 ;
        RECT 481.630 126.990 482.810 128.170 ;
        RECT 483.230 126.990 484.410 128.170 ;
        RECT 481.630 -26.910 482.810 -25.730 ;
        RECT 483.230 -26.910 484.410 -25.730 ;
        RECT 481.630 -28.510 482.810 -27.330 ;
        RECT 483.230 -28.510 484.410 -27.330 ;
        RECT 661.630 488.590 662.810 489.770 ;
        RECT 663.230 488.590 664.410 489.770 ;
        RECT 661.630 486.990 662.810 488.170 ;
        RECT 663.230 486.990 664.410 488.170 ;
        RECT 661.630 308.590 662.810 309.770 ;
        RECT 663.230 308.590 664.410 309.770 ;
        RECT 661.630 306.990 662.810 308.170 ;
        RECT 663.230 306.990 664.410 308.170 ;
        RECT 661.630 128.590 662.810 129.770 ;
        RECT 663.230 128.590 664.410 129.770 ;
        RECT 661.630 126.990 662.810 128.170 ;
        RECT 663.230 126.990 664.410 128.170 ;
        RECT 661.630 -26.910 662.810 -25.730 ;
        RECT 663.230 -26.910 664.410 -25.730 ;
        RECT 661.630 -28.510 662.810 -27.330 ;
        RECT 663.230 -28.510 664.410 -27.330 ;
        RECT 841.630 488.590 842.810 489.770 ;
        RECT 843.230 488.590 844.410 489.770 ;
        RECT 841.630 486.990 842.810 488.170 ;
        RECT 843.230 486.990 844.410 488.170 ;
        RECT 841.630 308.590 842.810 309.770 ;
        RECT 843.230 308.590 844.410 309.770 ;
        RECT 841.630 306.990 842.810 308.170 ;
        RECT 843.230 306.990 844.410 308.170 ;
        RECT 841.630 128.590 842.810 129.770 ;
        RECT 843.230 128.590 844.410 129.770 ;
        RECT 841.630 126.990 842.810 128.170 ;
        RECT 843.230 126.990 844.410 128.170 ;
        RECT 841.630 -26.910 842.810 -25.730 ;
        RECT 843.230 -26.910 844.410 -25.730 ;
        RECT 841.630 -28.510 842.810 -27.330 ;
        RECT 843.230 -28.510 844.410 -27.330 ;
        RECT 1021.630 3547.010 1022.810 3548.190 ;
        RECT 1023.230 3547.010 1024.410 3548.190 ;
        RECT 1021.630 3545.410 1022.810 3546.590 ;
        RECT 1023.230 3545.410 1024.410 3546.590 ;
        RECT 1021.630 3368.590 1022.810 3369.770 ;
        RECT 1023.230 3368.590 1024.410 3369.770 ;
        RECT 1021.630 3366.990 1022.810 3368.170 ;
        RECT 1023.230 3366.990 1024.410 3368.170 ;
        RECT 1021.630 3188.590 1022.810 3189.770 ;
        RECT 1023.230 3188.590 1024.410 3189.770 ;
        RECT 1021.630 3186.990 1022.810 3188.170 ;
        RECT 1023.230 3186.990 1024.410 3188.170 ;
        RECT 1021.630 3008.590 1022.810 3009.770 ;
        RECT 1023.230 3008.590 1024.410 3009.770 ;
        RECT 1021.630 3006.990 1022.810 3008.170 ;
        RECT 1023.230 3006.990 1024.410 3008.170 ;
        RECT 1021.630 2828.590 1022.810 2829.770 ;
        RECT 1023.230 2828.590 1024.410 2829.770 ;
        RECT 1021.630 2826.990 1022.810 2828.170 ;
        RECT 1023.230 2826.990 1024.410 2828.170 ;
        RECT 1021.630 2648.590 1022.810 2649.770 ;
        RECT 1023.230 2648.590 1024.410 2649.770 ;
        RECT 1021.630 2646.990 1022.810 2648.170 ;
        RECT 1023.230 2646.990 1024.410 2648.170 ;
        RECT 1021.630 2468.590 1022.810 2469.770 ;
        RECT 1023.230 2468.590 1024.410 2469.770 ;
        RECT 1021.630 2466.990 1022.810 2468.170 ;
        RECT 1023.230 2466.990 1024.410 2468.170 ;
        RECT 1021.630 2288.590 1022.810 2289.770 ;
        RECT 1023.230 2288.590 1024.410 2289.770 ;
        RECT 1021.630 2286.990 1022.810 2288.170 ;
        RECT 1023.230 2286.990 1024.410 2288.170 ;
        RECT 1021.630 2108.590 1022.810 2109.770 ;
        RECT 1023.230 2108.590 1024.410 2109.770 ;
        RECT 1021.630 2106.990 1022.810 2108.170 ;
        RECT 1023.230 2106.990 1024.410 2108.170 ;
        RECT 1021.630 1928.590 1022.810 1929.770 ;
        RECT 1023.230 1928.590 1024.410 1929.770 ;
        RECT 1021.630 1926.990 1022.810 1928.170 ;
        RECT 1023.230 1926.990 1024.410 1928.170 ;
        RECT 1021.630 1748.590 1022.810 1749.770 ;
        RECT 1023.230 1748.590 1024.410 1749.770 ;
        RECT 1021.630 1746.990 1022.810 1748.170 ;
        RECT 1023.230 1746.990 1024.410 1748.170 ;
        RECT 1021.630 1568.590 1022.810 1569.770 ;
        RECT 1023.230 1568.590 1024.410 1569.770 ;
        RECT 1021.630 1566.990 1022.810 1568.170 ;
        RECT 1023.230 1566.990 1024.410 1568.170 ;
        RECT 1021.630 1388.590 1022.810 1389.770 ;
        RECT 1023.230 1388.590 1024.410 1389.770 ;
        RECT 1021.630 1386.990 1022.810 1388.170 ;
        RECT 1023.230 1386.990 1024.410 1388.170 ;
        RECT 1021.630 1208.590 1022.810 1209.770 ;
        RECT 1023.230 1208.590 1024.410 1209.770 ;
        RECT 1021.630 1206.990 1022.810 1208.170 ;
        RECT 1023.230 1206.990 1024.410 1208.170 ;
        RECT 1021.630 1028.590 1022.810 1029.770 ;
        RECT 1023.230 1028.590 1024.410 1029.770 ;
        RECT 1021.630 1026.990 1022.810 1028.170 ;
        RECT 1023.230 1026.990 1024.410 1028.170 ;
        RECT 1021.630 848.590 1022.810 849.770 ;
        RECT 1023.230 848.590 1024.410 849.770 ;
        RECT 1021.630 846.990 1022.810 848.170 ;
        RECT 1023.230 846.990 1024.410 848.170 ;
        RECT 1021.630 668.590 1022.810 669.770 ;
        RECT 1023.230 668.590 1024.410 669.770 ;
        RECT 1021.630 666.990 1022.810 668.170 ;
        RECT 1023.230 666.990 1024.410 668.170 ;
        RECT 1021.630 488.590 1022.810 489.770 ;
        RECT 1023.230 488.590 1024.410 489.770 ;
        RECT 1021.630 486.990 1022.810 488.170 ;
        RECT 1023.230 486.990 1024.410 488.170 ;
        RECT 1021.630 308.590 1022.810 309.770 ;
        RECT 1023.230 308.590 1024.410 309.770 ;
        RECT 1021.630 306.990 1022.810 308.170 ;
        RECT 1023.230 306.990 1024.410 308.170 ;
        RECT 1021.630 128.590 1022.810 129.770 ;
        RECT 1023.230 128.590 1024.410 129.770 ;
        RECT 1021.630 126.990 1022.810 128.170 ;
        RECT 1023.230 126.990 1024.410 128.170 ;
        RECT 1021.630 -26.910 1022.810 -25.730 ;
        RECT 1023.230 -26.910 1024.410 -25.730 ;
        RECT 1021.630 -28.510 1022.810 -27.330 ;
        RECT 1023.230 -28.510 1024.410 -27.330 ;
        RECT 1201.630 3547.010 1202.810 3548.190 ;
        RECT 1203.230 3547.010 1204.410 3548.190 ;
        RECT 1201.630 3545.410 1202.810 3546.590 ;
        RECT 1203.230 3545.410 1204.410 3546.590 ;
        RECT 1201.630 3368.590 1202.810 3369.770 ;
        RECT 1203.230 3368.590 1204.410 3369.770 ;
        RECT 1201.630 3366.990 1202.810 3368.170 ;
        RECT 1203.230 3366.990 1204.410 3368.170 ;
        RECT 1201.630 3188.590 1202.810 3189.770 ;
        RECT 1203.230 3188.590 1204.410 3189.770 ;
        RECT 1201.630 3186.990 1202.810 3188.170 ;
        RECT 1203.230 3186.990 1204.410 3188.170 ;
        RECT 1201.630 3008.590 1202.810 3009.770 ;
        RECT 1203.230 3008.590 1204.410 3009.770 ;
        RECT 1201.630 3006.990 1202.810 3008.170 ;
        RECT 1203.230 3006.990 1204.410 3008.170 ;
        RECT 1201.630 2828.590 1202.810 2829.770 ;
        RECT 1203.230 2828.590 1204.410 2829.770 ;
        RECT 1201.630 2826.990 1202.810 2828.170 ;
        RECT 1203.230 2826.990 1204.410 2828.170 ;
        RECT 1201.630 2648.590 1202.810 2649.770 ;
        RECT 1203.230 2648.590 1204.410 2649.770 ;
        RECT 1201.630 2646.990 1202.810 2648.170 ;
        RECT 1203.230 2646.990 1204.410 2648.170 ;
        RECT 1201.630 2468.590 1202.810 2469.770 ;
        RECT 1203.230 2468.590 1204.410 2469.770 ;
        RECT 1201.630 2466.990 1202.810 2468.170 ;
        RECT 1203.230 2466.990 1204.410 2468.170 ;
        RECT 1201.630 2288.590 1202.810 2289.770 ;
        RECT 1203.230 2288.590 1204.410 2289.770 ;
        RECT 1201.630 2286.990 1202.810 2288.170 ;
        RECT 1203.230 2286.990 1204.410 2288.170 ;
        RECT 1201.630 2108.590 1202.810 2109.770 ;
        RECT 1203.230 2108.590 1204.410 2109.770 ;
        RECT 1201.630 2106.990 1202.810 2108.170 ;
        RECT 1203.230 2106.990 1204.410 2108.170 ;
        RECT 1201.630 1928.590 1202.810 1929.770 ;
        RECT 1203.230 1928.590 1204.410 1929.770 ;
        RECT 1201.630 1926.990 1202.810 1928.170 ;
        RECT 1203.230 1926.990 1204.410 1928.170 ;
        RECT 1201.630 1748.590 1202.810 1749.770 ;
        RECT 1203.230 1748.590 1204.410 1749.770 ;
        RECT 1201.630 1746.990 1202.810 1748.170 ;
        RECT 1203.230 1746.990 1204.410 1748.170 ;
        RECT 1201.630 1568.590 1202.810 1569.770 ;
        RECT 1203.230 1568.590 1204.410 1569.770 ;
        RECT 1201.630 1566.990 1202.810 1568.170 ;
        RECT 1203.230 1566.990 1204.410 1568.170 ;
        RECT 1201.630 1388.590 1202.810 1389.770 ;
        RECT 1203.230 1388.590 1204.410 1389.770 ;
        RECT 1201.630 1386.990 1202.810 1388.170 ;
        RECT 1203.230 1386.990 1204.410 1388.170 ;
        RECT 1201.630 1208.590 1202.810 1209.770 ;
        RECT 1203.230 1208.590 1204.410 1209.770 ;
        RECT 1201.630 1206.990 1202.810 1208.170 ;
        RECT 1203.230 1206.990 1204.410 1208.170 ;
        RECT 1201.630 1028.590 1202.810 1029.770 ;
        RECT 1203.230 1028.590 1204.410 1029.770 ;
        RECT 1201.630 1026.990 1202.810 1028.170 ;
        RECT 1203.230 1026.990 1204.410 1028.170 ;
        RECT 1201.630 848.590 1202.810 849.770 ;
        RECT 1203.230 848.590 1204.410 849.770 ;
        RECT 1201.630 846.990 1202.810 848.170 ;
        RECT 1203.230 846.990 1204.410 848.170 ;
        RECT 1201.630 668.590 1202.810 669.770 ;
        RECT 1203.230 668.590 1204.410 669.770 ;
        RECT 1201.630 666.990 1202.810 668.170 ;
        RECT 1203.230 666.990 1204.410 668.170 ;
        RECT 1201.630 488.590 1202.810 489.770 ;
        RECT 1203.230 488.590 1204.410 489.770 ;
        RECT 1201.630 486.990 1202.810 488.170 ;
        RECT 1203.230 486.990 1204.410 488.170 ;
        RECT 1201.630 308.590 1202.810 309.770 ;
        RECT 1203.230 308.590 1204.410 309.770 ;
        RECT 1201.630 306.990 1202.810 308.170 ;
        RECT 1203.230 306.990 1204.410 308.170 ;
        RECT 1201.630 128.590 1202.810 129.770 ;
        RECT 1203.230 128.590 1204.410 129.770 ;
        RECT 1201.630 126.990 1202.810 128.170 ;
        RECT 1203.230 126.990 1204.410 128.170 ;
        RECT 1201.630 -26.910 1202.810 -25.730 ;
        RECT 1203.230 -26.910 1204.410 -25.730 ;
        RECT 1201.630 -28.510 1202.810 -27.330 ;
        RECT 1203.230 -28.510 1204.410 -27.330 ;
        RECT 1381.630 3547.010 1382.810 3548.190 ;
        RECT 1383.230 3547.010 1384.410 3548.190 ;
        RECT 1381.630 3545.410 1382.810 3546.590 ;
        RECT 1383.230 3545.410 1384.410 3546.590 ;
        RECT 1381.630 3368.590 1382.810 3369.770 ;
        RECT 1383.230 3368.590 1384.410 3369.770 ;
        RECT 1381.630 3366.990 1382.810 3368.170 ;
        RECT 1383.230 3366.990 1384.410 3368.170 ;
        RECT 1381.630 3188.590 1382.810 3189.770 ;
        RECT 1383.230 3188.590 1384.410 3189.770 ;
        RECT 1381.630 3186.990 1382.810 3188.170 ;
        RECT 1383.230 3186.990 1384.410 3188.170 ;
        RECT 1381.630 3008.590 1382.810 3009.770 ;
        RECT 1383.230 3008.590 1384.410 3009.770 ;
        RECT 1381.630 3006.990 1382.810 3008.170 ;
        RECT 1383.230 3006.990 1384.410 3008.170 ;
        RECT 1381.630 2828.590 1382.810 2829.770 ;
        RECT 1383.230 2828.590 1384.410 2829.770 ;
        RECT 1381.630 2826.990 1382.810 2828.170 ;
        RECT 1383.230 2826.990 1384.410 2828.170 ;
        RECT 1381.630 2648.590 1382.810 2649.770 ;
        RECT 1383.230 2648.590 1384.410 2649.770 ;
        RECT 1381.630 2646.990 1382.810 2648.170 ;
        RECT 1383.230 2646.990 1384.410 2648.170 ;
        RECT 1381.630 2468.590 1382.810 2469.770 ;
        RECT 1383.230 2468.590 1384.410 2469.770 ;
        RECT 1381.630 2466.990 1382.810 2468.170 ;
        RECT 1383.230 2466.990 1384.410 2468.170 ;
        RECT 1381.630 2288.590 1382.810 2289.770 ;
        RECT 1383.230 2288.590 1384.410 2289.770 ;
        RECT 1381.630 2286.990 1382.810 2288.170 ;
        RECT 1383.230 2286.990 1384.410 2288.170 ;
        RECT 1381.630 2108.590 1382.810 2109.770 ;
        RECT 1383.230 2108.590 1384.410 2109.770 ;
        RECT 1381.630 2106.990 1382.810 2108.170 ;
        RECT 1383.230 2106.990 1384.410 2108.170 ;
        RECT 1381.630 1928.590 1382.810 1929.770 ;
        RECT 1383.230 1928.590 1384.410 1929.770 ;
        RECT 1381.630 1926.990 1382.810 1928.170 ;
        RECT 1383.230 1926.990 1384.410 1928.170 ;
        RECT 1381.630 1748.590 1382.810 1749.770 ;
        RECT 1383.230 1748.590 1384.410 1749.770 ;
        RECT 1381.630 1746.990 1382.810 1748.170 ;
        RECT 1383.230 1746.990 1384.410 1748.170 ;
        RECT 1381.630 1568.590 1382.810 1569.770 ;
        RECT 1383.230 1568.590 1384.410 1569.770 ;
        RECT 1381.630 1566.990 1382.810 1568.170 ;
        RECT 1383.230 1566.990 1384.410 1568.170 ;
        RECT 1381.630 1388.590 1382.810 1389.770 ;
        RECT 1383.230 1388.590 1384.410 1389.770 ;
        RECT 1381.630 1386.990 1382.810 1388.170 ;
        RECT 1383.230 1386.990 1384.410 1388.170 ;
        RECT 1381.630 1208.590 1382.810 1209.770 ;
        RECT 1383.230 1208.590 1384.410 1209.770 ;
        RECT 1381.630 1206.990 1382.810 1208.170 ;
        RECT 1383.230 1206.990 1384.410 1208.170 ;
        RECT 1381.630 1028.590 1382.810 1029.770 ;
        RECT 1383.230 1028.590 1384.410 1029.770 ;
        RECT 1381.630 1026.990 1382.810 1028.170 ;
        RECT 1383.230 1026.990 1384.410 1028.170 ;
        RECT 1381.630 848.590 1382.810 849.770 ;
        RECT 1383.230 848.590 1384.410 849.770 ;
        RECT 1381.630 846.990 1382.810 848.170 ;
        RECT 1383.230 846.990 1384.410 848.170 ;
        RECT 1381.630 668.590 1382.810 669.770 ;
        RECT 1383.230 668.590 1384.410 669.770 ;
        RECT 1381.630 666.990 1382.810 668.170 ;
        RECT 1383.230 666.990 1384.410 668.170 ;
        RECT 1381.630 488.590 1382.810 489.770 ;
        RECT 1383.230 488.590 1384.410 489.770 ;
        RECT 1381.630 486.990 1382.810 488.170 ;
        RECT 1383.230 486.990 1384.410 488.170 ;
        RECT 1381.630 308.590 1382.810 309.770 ;
        RECT 1383.230 308.590 1384.410 309.770 ;
        RECT 1381.630 306.990 1382.810 308.170 ;
        RECT 1383.230 306.990 1384.410 308.170 ;
        RECT 1381.630 128.590 1382.810 129.770 ;
        RECT 1383.230 128.590 1384.410 129.770 ;
        RECT 1381.630 126.990 1382.810 128.170 ;
        RECT 1383.230 126.990 1384.410 128.170 ;
        RECT 1381.630 -26.910 1382.810 -25.730 ;
        RECT 1383.230 -26.910 1384.410 -25.730 ;
        RECT 1381.630 -28.510 1382.810 -27.330 ;
        RECT 1383.230 -28.510 1384.410 -27.330 ;
        RECT 1561.630 3547.010 1562.810 3548.190 ;
        RECT 1563.230 3547.010 1564.410 3548.190 ;
        RECT 1561.630 3545.410 1562.810 3546.590 ;
        RECT 1563.230 3545.410 1564.410 3546.590 ;
        RECT 1561.630 3368.590 1562.810 3369.770 ;
        RECT 1563.230 3368.590 1564.410 3369.770 ;
        RECT 1561.630 3366.990 1562.810 3368.170 ;
        RECT 1563.230 3366.990 1564.410 3368.170 ;
        RECT 1561.630 3188.590 1562.810 3189.770 ;
        RECT 1563.230 3188.590 1564.410 3189.770 ;
        RECT 1561.630 3186.990 1562.810 3188.170 ;
        RECT 1563.230 3186.990 1564.410 3188.170 ;
        RECT 1561.630 3008.590 1562.810 3009.770 ;
        RECT 1563.230 3008.590 1564.410 3009.770 ;
        RECT 1561.630 3006.990 1562.810 3008.170 ;
        RECT 1563.230 3006.990 1564.410 3008.170 ;
        RECT 1561.630 2828.590 1562.810 2829.770 ;
        RECT 1563.230 2828.590 1564.410 2829.770 ;
        RECT 1561.630 2826.990 1562.810 2828.170 ;
        RECT 1563.230 2826.990 1564.410 2828.170 ;
        RECT 1561.630 2648.590 1562.810 2649.770 ;
        RECT 1563.230 2648.590 1564.410 2649.770 ;
        RECT 1561.630 2646.990 1562.810 2648.170 ;
        RECT 1563.230 2646.990 1564.410 2648.170 ;
        RECT 1561.630 2468.590 1562.810 2469.770 ;
        RECT 1563.230 2468.590 1564.410 2469.770 ;
        RECT 1561.630 2466.990 1562.810 2468.170 ;
        RECT 1563.230 2466.990 1564.410 2468.170 ;
        RECT 1561.630 2288.590 1562.810 2289.770 ;
        RECT 1563.230 2288.590 1564.410 2289.770 ;
        RECT 1561.630 2286.990 1562.810 2288.170 ;
        RECT 1563.230 2286.990 1564.410 2288.170 ;
        RECT 1561.630 2108.590 1562.810 2109.770 ;
        RECT 1563.230 2108.590 1564.410 2109.770 ;
        RECT 1561.630 2106.990 1562.810 2108.170 ;
        RECT 1563.230 2106.990 1564.410 2108.170 ;
        RECT 1561.630 1928.590 1562.810 1929.770 ;
        RECT 1563.230 1928.590 1564.410 1929.770 ;
        RECT 1561.630 1926.990 1562.810 1928.170 ;
        RECT 1563.230 1926.990 1564.410 1928.170 ;
        RECT 1561.630 1748.590 1562.810 1749.770 ;
        RECT 1563.230 1748.590 1564.410 1749.770 ;
        RECT 1561.630 1746.990 1562.810 1748.170 ;
        RECT 1563.230 1746.990 1564.410 1748.170 ;
        RECT 1561.630 1568.590 1562.810 1569.770 ;
        RECT 1563.230 1568.590 1564.410 1569.770 ;
        RECT 1561.630 1566.990 1562.810 1568.170 ;
        RECT 1563.230 1566.990 1564.410 1568.170 ;
        RECT 1561.630 1388.590 1562.810 1389.770 ;
        RECT 1563.230 1388.590 1564.410 1389.770 ;
        RECT 1561.630 1386.990 1562.810 1388.170 ;
        RECT 1563.230 1386.990 1564.410 1388.170 ;
        RECT 1561.630 1208.590 1562.810 1209.770 ;
        RECT 1563.230 1208.590 1564.410 1209.770 ;
        RECT 1561.630 1206.990 1562.810 1208.170 ;
        RECT 1563.230 1206.990 1564.410 1208.170 ;
        RECT 1561.630 1028.590 1562.810 1029.770 ;
        RECT 1563.230 1028.590 1564.410 1029.770 ;
        RECT 1561.630 1026.990 1562.810 1028.170 ;
        RECT 1563.230 1026.990 1564.410 1028.170 ;
        RECT 1561.630 848.590 1562.810 849.770 ;
        RECT 1563.230 848.590 1564.410 849.770 ;
        RECT 1561.630 846.990 1562.810 848.170 ;
        RECT 1563.230 846.990 1564.410 848.170 ;
        RECT 1561.630 668.590 1562.810 669.770 ;
        RECT 1563.230 668.590 1564.410 669.770 ;
        RECT 1561.630 666.990 1562.810 668.170 ;
        RECT 1563.230 666.990 1564.410 668.170 ;
        RECT 1561.630 488.590 1562.810 489.770 ;
        RECT 1563.230 488.590 1564.410 489.770 ;
        RECT 1561.630 486.990 1562.810 488.170 ;
        RECT 1563.230 486.990 1564.410 488.170 ;
        RECT 1561.630 308.590 1562.810 309.770 ;
        RECT 1563.230 308.590 1564.410 309.770 ;
        RECT 1561.630 306.990 1562.810 308.170 ;
        RECT 1563.230 306.990 1564.410 308.170 ;
        RECT 1561.630 128.590 1562.810 129.770 ;
        RECT 1563.230 128.590 1564.410 129.770 ;
        RECT 1561.630 126.990 1562.810 128.170 ;
        RECT 1563.230 126.990 1564.410 128.170 ;
        RECT 1561.630 -26.910 1562.810 -25.730 ;
        RECT 1563.230 -26.910 1564.410 -25.730 ;
        RECT 1561.630 -28.510 1562.810 -27.330 ;
        RECT 1563.230 -28.510 1564.410 -27.330 ;
        RECT 1741.630 3547.010 1742.810 3548.190 ;
        RECT 1743.230 3547.010 1744.410 3548.190 ;
        RECT 1741.630 3545.410 1742.810 3546.590 ;
        RECT 1743.230 3545.410 1744.410 3546.590 ;
        RECT 1741.630 3368.590 1742.810 3369.770 ;
        RECT 1743.230 3368.590 1744.410 3369.770 ;
        RECT 1741.630 3366.990 1742.810 3368.170 ;
        RECT 1743.230 3366.990 1744.410 3368.170 ;
        RECT 1741.630 3188.590 1742.810 3189.770 ;
        RECT 1743.230 3188.590 1744.410 3189.770 ;
        RECT 1741.630 3186.990 1742.810 3188.170 ;
        RECT 1743.230 3186.990 1744.410 3188.170 ;
        RECT 1741.630 3008.590 1742.810 3009.770 ;
        RECT 1743.230 3008.590 1744.410 3009.770 ;
        RECT 1741.630 3006.990 1742.810 3008.170 ;
        RECT 1743.230 3006.990 1744.410 3008.170 ;
        RECT 1741.630 2828.590 1742.810 2829.770 ;
        RECT 1743.230 2828.590 1744.410 2829.770 ;
        RECT 1741.630 2826.990 1742.810 2828.170 ;
        RECT 1743.230 2826.990 1744.410 2828.170 ;
        RECT 1741.630 2648.590 1742.810 2649.770 ;
        RECT 1743.230 2648.590 1744.410 2649.770 ;
        RECT 1741.630 2646.990 1742.810 2648.170 ;
        RECT 1743.230 2646.990 1744.410 2648.170 ;
        RECT 1741.630 2468.590 1742.810 2469.770 ;
        RECT 1743.230 2468.590 1744.410 2469.770 ;
        RECT 1741.630 2466.990 1742.810 2468.170 ;
        RECT 1743.230 2466.990 1744.410 2468.170 ;
        RECT 1741.630 2288.590 1742.810 2289.770 ;
        RECT 1743.230 2288.590 1744.410 2289.770 ;
        RECT 1741.630 2286.990 1742.810 2288.170 ;
        RECT 1743.230 2286.990 1744.410 2288.170 ;
        RECT 1741.630 2108.590 1742.810 2109.770 ;
        RECT 1743.230 2108.590 1744.410 2109.770 ;
        RECT 1741.630 2106.990 1742.810 2108.170 ;
        RECT 1743.230 2106.990 1744.410 2108.170 ;
        RECT 1741.630 1928.590 1742.810 1929.770 ;
        RECT 1743.230 1928.590 1744.410 1929.770 ;
        RECT 1741.630 1926.990 1742.810 1928.170 ;
        RECT 1743.230 1926.990 1744.410 1928.170 ;
        RECT 1741.630 1748.590 1742.810 1749.770 ;
        RECT 1743.230 1748.590 1744.410 1749.770 ;
        RECT 1741.630 1746.990 1742.810 1748.170 ;
        RECT 1743.230 1746.990 1744.410 1748.170 ;
        RECT 1741.630 1568.590 1742.810 1569.770 ;
        RECT 1743.230 1568.590 1744.410 1569.770 ;
        RECT 1741.630 1566.990 1742.810 1568.170 ;
        RECT 1743.230 1566.990 1744.410 1568.170 ;
        RECT 1741.630 1388.590 1742.810 1389.770 ;
        RECT 1743.230 1388.590 1744.410 1389.770 ;
        RECT 1741.630 1386.990 1742.810 1388.170 ;
        RECT 1743.230 1386.990 1744.410 1388.170 ;
        RECT 1741.630 1208.590 1742.810 1209.770 ;
        RECT 1743.230 1208.590 1744.410 1209.770 ;
        RECT 1741.630 1206.990 1742.810 1208.170 ;
        RECT 1743.230 1206.990 1744.410 1208.170 ;
        RECT 1741.630 1028.590 1742.810 1029.770 ;
        RECT 1743.230 1028.590 1744.410 1029.770 ;
        RECT 1741.630 1026.990 1742.810 1028.170 ;
        RECT 1743.230 1026.990 1744.410 1028.170 ;
        RECT 1741.630 848.590 1742.810 849.770 ;
        RECT 1743.230 848.590 1744.410 849.770 ;
        RECT 1741.630 846.990 1742.810 848.170 ;
        RECT 1743.230 846.990 1744.410 848.170 ;
        RECT 1741.630 668.590 1742.810 669.770 ;
        RECT 1743.230 668.590 1744.410 669.770 ;
        RECT 1741.630 666.990 1742.810 668.170 ;
        RECT 1743.230 666.990 1744.410 668.170 ;
        RECT 1741.630 488.590 1742.810 489.770 ;
        RECT 1743.230 488.590 1744.410 489.770 ;
        RECT 1741.630 486.990 1742.810 488.170 ;
        RECT 1743.230 486.990 1744.410 488.170 ;
        RECT 1741.630 308.590 1742.810 309.770 ;
        RECT 1743.230 308.590 1744.410 309.770 ;
        RECT 1741.630 306.990 1742.810 308.170 ;
        RECT 1743.230 306.990 1744.410 308.170 ;
        RECT 1741.630 128.590 1742.810 129.770 ;
        RECT 1743.230 128.590 1744.410 129.770 ;
        RECT 1741.630 126.990 1742.810 128.170 ;
        RECT 1743.230 126.990 1744.410 128.170 ;
        RECT 1741.630 -26.910 1742.810 -25.730 ;
        RECT 1743.230 -26.910 1744.410 -25.730 ;
        RECT 1741.630 -28.510 1742.810 -27.330 ;
        RECT 1743.230 -28.510 1744.410 -27.330 ;
        RECT 1921.630 3547.010 1922.810 3548.190 ;
        RECT 1923.230 3547.010 1924.410 3548.190 ;
        RECT 1921.630 3545.410 1922.810 3546.590 ;
        RECT 1923.230 3545.410 1924.410 3546.590 ;
        RECT 1921.630 3368.590 1922.810 3369.770 ;
        RECT 1923.230 3368.590 1924.410 3369.770 ;
        RECT 1921.630 3366.990 1922.810 3368.170 ;
        RECT 1923.230 3366.990 1924.410 3368.170 ;
        RECT 1921.630 3188.590 1922.810 3189.770 ;
        RECT 1923.230 3188.590 1924.410 3189.770 ;
        RECT 1921.630 3186.990 1922.810 3188.170 ;
        RECT 1923.230 3186.990 1924.410 3188.170 ;
        RECT 1921.630 3008.590 1922.810 3009.770 ;
        RECT 1923.230 3008.590 1924.410 3009.770 ;
        RECT 1921.630 3006.990 1922.810 3008.170 ;
        RECT 1923.230 3006.990 1924.410 3008.170 ;
        RECT 1921.630 2828.590 1922.810 2829.770 ;
        RECT 1923.230 2828.590 1924.410 2829.770 ;
        RECT 1921.630 2826.990 1922.810 2828.170 ;
        RECT 1923.230 2826.990 1924.410 2828.170 ;
        RECT 1921.630 2648.590 1922.810 2649.770 ;
        RECT 1923.230 2648.590 1924.410 2649.770 ;
        RECT 1921.630 2646.990 1922.810 2648.170 ;
        RECT 1923.230 2646.990 1924.410 2648.170 ;
        RECT 1921.630 2468.590 1922.810 2469.770 ;
        RECT 1923.230 2468.590 1924.410 2469.770 ;
        RECT 1921.630 2466.990 1922.810 2468.170 ;
        RECT 1923.230 2466.990 1924.410 2468.170 ;
        RECT 1921.630 2288.590 1922.810 2289.770 ;
        RECT 1923.230 2288.590 1924.410 2289.770 ;
        RECT 1921.630 2286.990 1922.810 2288.170 ;
        RECT 1923.230 2286.990 1924.410 2288.170 ;
        RECT 1921.630 2108.590 1922.810 2109.770 ;
        RECT 1923.230 2108.590 1924.410 2109.770 ;
        RECT 1921.630 2106.990 1922.810 2108.170 ;
        RECT 1923.230 2106.990 1924.410 2108.170 ;
        RECT 1921.630 1928.590 1922.810 1929.770 ;
        RECT 1923.230 1928.590 1924.410 1929.770 ;
        RECT 1921.630 1926.990 1922.810 1928.170 ;
        RECT 1923.230 1926.990 1924.410 1928.170 ;
        RECT 1921.630 1748.590 1922.810 1749.770 ;
        RECT 1923.230 1748.590 1924.410 1749.770 ;
        RECT 1921.630 1746.990 1922.810 1748.170 ;
        RECT 1923.230 1746.990 1924.410 1748.170 ;
        RECT 1921.630 1568.590 1922.810 1569.770 ;
        RECT 1923.230 1568.590 1924.410 1569.770 ;
        RECT 1921.630 1566.990 1922.810 1568.170 ;
        RECT 1923.230 1566.990 1924.410 1568.170 ;
        RECT 1921.630 1388.590 1922.810 1389.770 ;
        RECT 1923.230 1388.590 1924.410 1389.770 ;
        RECT 1921.630 1386.990 1922.810 1388.170 ;
        RECT 1923.230 1386.990 1924.410 1388.170 ;
        RECT 1921.630 1208.590 1922.810 1209.770 ;
        RECT 1923.230 1208.590 1924.410 1209.770 ;
        RECT 1921.630 1206.990 1922.810 1208.170 ;
        RECT 1923.230 1206.990 1924.410 1208.170 ;
        RECT 1921.630 1028.590 1922.810 1029.770 ;
        RECT 1923.230 1028.590 1924.410 1029.770 ;
        RECT 1921.630 1026.990 1922.810 1028.170 ;
        RECT 1923.230 1026.990 1924.410 1028.170 ;
        RECT 1921.630 848.590 1922.810 849.770 ;
        RECT 1923.230 848.590 1924.410 849.770 ;
        RECT 1921.630 846.990 1922.810 848.170 ;
        RECT 1923.230 846.990 1924.410 848.170 ;
        RECT 1921.630 668.590 1922.810 669.770 ;
        RECT 1923.230 668.590 1924.410 669.770 ;
        RECT 1921.630 666.990 1922.810 668.170 ;
        RECT 1923.230 666.990 1924.410 668.170 ;
        RECT 1921.630 488.590 1922.810 489.770 ;
        RECT 1923.230 488.590 1924.410 489.770 ;
        RECT 1921.630 486.990 1922.810 488.170 ;
        RECT 1923.230 486.990 1924.410 488.170 ;
        RECT 1921.630 308.590 1922.810 309.770 ;
        RECT 1923.230 308.590 1924.410 309.770 ;
        RECT 1921.630 306.990 1922.810 308.170 ;
        RECT 1923.230 306.990 1924.410 308.170 ;
        RECT 1921.630 128.590 1922.810 129.770 ;
        RECT 1923.230 128.590 1924.410 129.770 ;
        RECT 1921.630 126.990 1922.810 128.170 ;
        RECT 1923.230 126.990 1924.410 128.170 ;
        RECT 1921.630 -26.910 1922.810 -25.730 ;
        RECT 1923.230 -26.910 1924.410 -25.730 ;
        RECT 1921.630 -28.510 1922.810 -27.330 ;
        RECT 1923.230 -28.510 1924.410 -27.330 ;
        RECT 2101.630 3547.010 2102.810 3548.190 ;
        RECT 2103.230 3547.010 2104.410 3548.190 ;
        RECT 2101.630 3545.410 2102.810 3546.590 ;
        RECT 2103.230 3545.410 2104.410 3546.590 ;
        RECT 2101.630 3368.590 2102.810 3369.770 ;
        RECT 2103.230 3368.590 2104.410 3369.770 ;
        RECT 2101.630 3366.990 2102.810 3368.170 ;
        RECT 2103.230 3366.990 2104.410 3368.170 ;
        RECT 2101.630 3188.590 2102.810 3189.770 ;
        RECT 2103.230 3188.590 2104.410 3189.770 ;
        RECT 2101.630 3186.990 2102.810 3188.170 ;
        RECT 2103.230 3186.990 2104.410 3188.170 ;
        RECT 2101.630 3008.590 2102.810 3009.770 ;
        RECT 2103.230 3008.590 2104.410 3009.770 ;
        RECT 2101.630 3006.990 2102.810 3008.170 ;
        RECT 2103.230 3006.990 2104.410 3008.170 ;
        RECT 2101.630 2828.590 2102.810 2829.770 ;
        RECT 2103.230 2828.590 2104.410 2829.770 ;
        RECT 2101.630 2826.990 2102.810 2828.170 ;
        RECT 2103.230 2826.990 2104.410 2828.170 ;
        RECT 2101.630 2648.590 2102.810 2649.770 ;
        RECT 2103.230 2648.590 2104.410 2649.770 ;
        RECT 2101.630 2646.990 2102.810 2648.170 ;
        RECT 2103.230 2646.990 2104.410 2648.170 ;
        RECT 2101.630 2468.590 2102.810 2469.770 ;
        RECT 2103.230 2468.590 2104.410 2469.770 ;
        RECT 2101.630 2466.990 2102.810 2468.170 ;
        RECT 2103.230 2466.990 2104.410 2468.170 ;
        RECT 2101.630 2288.590 2102.810 2289.770 ;
        RECT 2103.230 2288.590 2104.410 2289.770 ;
        RECT 2101.630 2286.990 2102.810 2288.170 ;
        RECT 2103.230 2286.990 2104.410 2288.170 ;
        RECT 2101.630 2108.590 2102.810 2109.770 ;
        RECT 2103.230 2108.590 2104.410 2109.770 ;
        RECT 2101.630 2106.990 2102.810 2108.170 ;
        RECT 2103.230 2106.990 2104.410 2108.170 ;
        RECT 2101.630 1928.590 2102.810 1929.770 ;
        RECT 2103.230 1928.590 2104.410 1929.770 ;
        RECT 2101.630 1926.990 2102.810 1928.170 ;
        RECT 2103.230 1926.990 2104.410 1928.170 ;
        RECT 2101.630 1748.590 2102.810 1749.770 ;
        RECT 2103.230 1748.590 2104.410 1749.770 ;
        RECT 2101.630 1746.990 2102.810 1748.170 ;
        RECT 2103.230 1746.990 2104.410 1748.170 ;
        RECT 2101.630 1568.590 2102.810 1569.770 ;
        RECT 2103.230 1568.590 2104.410 1569.770 ;
        RECT 2101.630 1566.990 2102.810 1568.170 ;
        RECT 2103.230 1566.990 2104.410 1568.170 ;
        RECT 2101.630 1388.590 2102.810 1389.770 ;
        RECT 2103.230 1388.590 2104.410 1389.770 ;
        RECT 2101.630 1386.990 2102.810 1388.170 ;
        RECT 2103.230 1386.990 2104.410 1388.170 ;
        RECT 2101.630 1208.590 2102.810 1209.770 ;
        RECT 2103.230 1208.590 2104.410 1209.770 ;
        RECT 2101.630 1206.990 2102.810 1208.170 ;
        RECT 2103.230 1206.990 2104.410 1208.170 ;
        RECT 2101.630 1028.590 2102.810 1029.770 ;
        RECT 2103.230 1028.590 2104.410 1029.770 ;
        RECT 2101.630 1026.990 2102.810 1028.170 ;
        RECT 2103.230 1026.990 2104.410 1028.170 ;
        RECT 2101.630 848.590 2102.810 849.770 ;
        RECT 2103.230 848.590 2104.410 849.770 ;
        RECT 2101.630 846.990 2102.810 848.170 ;
        RECT 2103.230 846.990 2104.410 848.170 ;
        RECT 2101.630 668.590 2102.810 669.770 ;
        RECT 2103.230 668.590 2104.410 669.770 ;
        RECT 2101.630 666.990 2102.810 668.170 ;
        RECT 2103.230 666.990 2104.410 668.170 ;
        RECT 2101.630 488.590 2102.810 489.770 ;
        RECT 2103.230 488.590 2104.410 489.770 ;
        RECT 2101.630 486.990 2102.810 488.170 ;
        RECT 2103.230 486.990 2104.410 488.170 ;
        RECT 2101.630 308.590 2102.810 309.770 ;
        RECT 2103.230 308.590 2104.410 309.770 ;
        RECT 2101.630 306.990 2102.810 308.170 ;
        RECT 2103.230 306.990 2104.410 308.170 ;
        RECT 2101.630 128.590 2102.810 129.770 ;
        RECT 2103.230 128.590 2104.410 129.770 ;
        RECT 2101.630 126.990 2102.810 128.170 ;
        RECT 2103.230 126.990 2104.410 128.170 ;
        RECT 2101.630 -26.910 2102.810 -25.730 ;
        RECT 2103.230 -26.910 2104.410 -25.730 ;
        RECT 2101.630 -28.510 2102.810 -27.330 ;
        RECT 2103.230 -28.510 2104.410 -27.330 ;
        RECT 2281.630 3547.010 2282.810 3548.190 ;
        RECT 2283.230 3547.010 2284.410 3548.190 ;
        RECT 2281.630 3545.410 2282.810 3546.590 ;
        RECT 2283.230 3545.410 2284.410 3546.590 ;
        RECT 2281.630 3368.590 2282.810 3369.770 ;
        RECT 2283.230 3368.590 2284.410 3369.770 ;
        RECT 2281.630 3366.990 2282.810 3368.170 ;
        RECT 2283.230 3366.990 2284.410 3368.170 ;
        RECT 2281.630 3188.590 2282.810 3189.770 ;
        RECT 2283.230 3188.590 2284.410 3189.770 ;
        RECT 2281.630 3186.990 2282.810 3188.170 ;
        RECT 2283.230 3186.990 2284.410 3188.170 ;
        RECT 2281.630 3008.590 2282.810 3009.770 ;
        RECT 2283.230 3008.590 2284.410 3009.770 ;
        RECT 2281.630 3006.990 2282.810 3008.170 ;
        RECT 2283.230 3006.990 2284.410 3008.170 ;
        RECT 2281.630 2828.590 2282.810 2829.770 ;
        RECT 2283.230 2828.590 2284.410 2829.770 ;
        RECT 2281.630 2826.990 2282.810 2828.170 ;
        RECT 2283.230 2826.990 2284.410 2828.170 ;
        RECT 2281.630 2648.590 2282.810 2649.770 ;
        RECT 2283.230 2648.590 2284.410 2649.770 ;
        RECT 2281.630 2646.990 2282.810 2648.170 ;
        RECT 2283.230 2646.990 2284.410 2648.170 ;
        RECT 2281.630 2468.590 2282.810 2469.770 ;
        RECT 2283.230 2468.590 2284.410 2469.770 ;
        RECT 2281.630 2466.990 2282.810 2468.170 ;
        RECT 2283.230 2466.990 2284.410 2468.170 ;
        RECT 2281.630 2288.590 2282.810 2289.770 ;
        RECT 2283.230 2288.590 2284.410 2289.770 ;
        RECT 2281.630 2286.990 2282.810 2288.170 ;
        RECT 2283.230 2286.990 2284.410 2288.170 ;
        RECT 2281.630 2108.590 2282.810 2109.770 ;
        RECT 2283.230 2108.590 2284.410 2109.770 ;
        RECT 2281.630 2106.990 2282.810 2108.170 ;
        RECT 2283.230 2106.990 2284.410 2108.170 ;
        RECT 2281.630 1928.590 2282.810 1929.770 ;
        RECT 2283.230 1928.590 2284.410 1929.770 ;
        RECT 2281.630 1926.990 2282.810 1928.170 ;
        RECT 2283.230 1926.990 2284.410 1928.170 ;
        RECT 2281.630 1748.590 2282.810 1749.770 ;
        RECT 2283.230 1748.590 2284.410 1749.770 ;
        RECT 2281.630 1746.990 2282.810 1748.170 ;
        RECT 2283.230 1746.990 2284.410 1748.170 ;
        RECT 2281.630 1568.590 2282.810 1569.770 ;
        RECT 2283.230 1568.590 2284.410 1569.770 ;
        RECT 2281.630 1566.990 2282.810 1568.170 ;
        RECT 2283.230 1566.990 2284.410 1568.170 ;
        RECT 2281.630 1388.590 2282.810 1389.770 ;
        RECT 2283.230 1388.590 2284.410 1389.770 ;
        RECT 2281.630 1386.990 2282.810 1388.170 ;
        RECT 2283.230 1386.990 2284.410 1388.170 ;
        RECT 2281.630 1208.590 2282.810 1209.770 ;
        RECT 2283.230 1208.590 2284.410 1209.770 ;
        RECT 2281.630 1206.990 2282.810 1208.170 ;
        RECT 2283.230 1206.990 2284.410 1208.170 ;
        RECT 2281.630 1028.590 2282.810 1029.770 ;
        RECT 2283.230 1028.590 2284.410 1029.770 ;
        RECT 2281.630 1026.990 2282.810 1028.170 ;
        RECT 2283.230 1026.990 2284.410 1028.170 ;
        RECT 2281.630 848.590 2282.810 849.770 ;
        RECT 2283.230 848.590 2284.410 849.770 ;
        RECT 2281.630 846.990 2282.810 848.170 ;
        RECT 2283.230 846.990 2284.410 848.170 ;
        RECT 2281.630 668.590 2282.810 669.770 ;
        RECT 2283.230 668.590 2284.410 669.770 ;
        RECT 2281.630 666.990 2282.810 668.170 ;
        RECT 2283.230 666.990 2284.410 668.170 ;
        RECT 2281.630 488.590 2282.810 489.770 ;
        RECT 2283.230 488.590 2284.410 489.770 ;
        RECT 2281.630 486.990 2282.810 488.170 ;
        RECT 2283.230 486.990 2284.410 488.170 ;
        RECT 2281.630 308.590 2282.810 309.770 ;
        RECT 2283.230 308.590 2284.410 309.770 ;
        RECT 2281.630 306.990 2282.810 308.170 ;
        RECT 2283.230 306.990 2284.410 308.170 ;
        RECT 2281.630 128.590 2282.810 129.770 ;
        RECT 2283.230 128.590 2284.410 129.770 ;
        RECT 2281.630 126.990 2282.810 128.170 ;
        RECT 2283.230 126.990 2284.410 128.170 ;
        RECT 2281.630 -26.910 2282.810 -25.730 ;
        RECT 2283.230 -26.910 2284.410 -25.730 ;
        RECT 2281.630 -28.510 2282.810 -27.330 ;
        RECT 2283.230 -28.510 2284.410 -27.330 ;
        RECT 2461.630 3547.010 2462.810 3548.190 ;
        RECT 2463.230 3547.010 2464.410 3548.190 ;
        RECT 2461.630 3545.410 2462.810 3546.590 ;
        RECT 2463.230 3545.410 2464.410 3546.590 ;
        RECT 2461.630 3368.590 2462.810 3369.770 ;
        RECT 2463.230 3368.590 2464.410 3369.770 ;
        RECT 2461.630 3366.990 2462.810 3368.170 ;
        RECT 2463.230 3366.990 2464.410 3368.170 ;
        RECT 2461.630 3188.590 2462.810 3189.770 ;
        RECT 2463.230 3188.590 2464.410 3189.770 ;
        RECT 2461.630 3186.990 2462.810 3188.170 ;
        RECT 2463.230 3186.990 2464.410 3188.170 ;
        RECT 2461.630 3008.590 2462.810 3009.770 ;
        RECT 2463.230 3008.590 2464.410 3009.770 ;
        RECT 2461.630 3006.990 2462.810 3008.170 ;
        RECT 2463.230 3006.990 2464.410 3008.170 ;
        RECT 2461.630 2828.590 2462.810 2829.770 ;
        RECT 2463.230 2828.590 2464.410 2829.770 ;
        RECT 2461.630 2826.990 2462.810 2828.170 ;
        RECT 2463.230 2826.990 2464.410 2828.170 ;
        RECT 2461.630 2648.590 2462.810 2649.770 ;
        RECT 2463.230 2648.590 2464.410 2649.770 ;
        RECT 2461.630 2646.990 2462.810 2648.170 ;
        RECT 2463.230 2646.990 2464.410 2648.170 ;
        RECT 2461.630 2468.590 2462.810 2469.770 ;
        RECT 2463.230 2468.590 2464.410 2469.770 ;
        RECT 2461.630 2466.990 2462.810 2468.170 ;
        RECT 2463.230 2466.990 2464.410 2468.170 ;
        RECT 2461.630 2288.590 2462.810 2289.770 ;
        RECT 2463.230 2288.590 2464.410 2289.770 ;
        RECT 2461.630 2286.990 2462.810 2288.170 ;
        RECT 2463.230 2286.990 2464.410 2288.170 ;
        RECT 2461.630 2108.590 2462.810 2109.770 ;
        RECT 2463.230 2108.590 2464.410 2109.770 ;
        RECT 2461.630 2106.990 2462.810 2108.170 ;
        RECT 2463.230 2106.990 2464.410 2108.170 ;
        RECT 2461.630 1928.590 2462.810 1929.770 ;
        RECT 2463.230 1928.590 2464.410 1929.770 ;
        RECT 2461.630 1926.990 2462.810 1928.170 ;
        RECT 2463.230 1926.990 2464.410 1928.170 ;
        RECT 2461.630 1748.590 2462.810 1749.770 ;
        RECT 2463.230 1748.590 2464.410 1749.770 ;
        RECT 2461.630 1746.990 2462.810 1748.170 ;
        RECT 2463.230 1746.990 2464.410 1748.170 ;
        RECT 2461.630 1568.590 2462.810 1569.770 ;
        RECT 2463.230 1568.590 2464.410 1569.770 ;
        RECT 2461.630 1566.990 2462.810 1568.170 ;
        RECT 2463.230 1566.990 2464.410 1568.170 ;
        RECT 2461.630 1388.590 2462.810 1389.770 ;
        RECT 2463.230 1388.590 2464.410 1389.770 ;
        RECT 2461.630 1386.990 2462.810 1388.170 ;
        RECT 2463.230 1386.990 2464.410 1388.170 ;
        RECT 2461.630 1208.590 2462.810 1209.770 ;
        RECT 2463.230 1208.590 2464.410 1209.770 ;
        RECT 2461.630 1206.990 2462.810 1208.170 ;
        RECT 2463.230 1206.990 2464.410 1208.170 ;
        RECT 2461.630 1028.590 2462.810 1029.770 ;
        RECT 2463.230 1028.590 2464.410 1029.770 ;
        RECT 2461.630 1026.990 2462.810 1028.170 ;
        RECT 2463.230 1026.990 2464.410 1028.170 ;
        RECT 2461.630 848.590 2462.810 849.770 ;
        RECT 2463.230 848.590 2464.410 849.770 ;
        RECT 2461.630 846.990 2462.810 848.170 ;
        RECT 2463.230 846.990 2464.410 848.170 ;
        RECT 2461.630 668.590 2462.810 669.770 ;
        RECT 2463.230 668.590 2464.410 669.770 ;
        RECT 2461.630 666.990 2462.810 668.170 ;
        RECT 2463.230 666.990 2464.410 668.170 ;
        RECT 2461.630 488.590 2462.810 489.770 ;
        RECT 2463.230 488.590 2464.410 489.770 ;
        RECT 2461.630 486.990 2462.810 488.170 ;
        RECT 2463.230 486.990 2464.410 488.170 ;
        RECT 2461.630 308.590 2462.810 309.770 ;
        RECT 2463.230 308.590 2464.410 309.770 ;
        RECT 2461.630 306.990 2462.810 308.170 ;
        RECT 2463.230 306.990 2464.410 308.170 ;
        RECT 2461.630 128.590 2462.810 129.770 ;
        RECT 2463.230 128.590 2464.410 129.770 ;
        RECT 2461.630 126.990 2462.810 128.170 ;
        RECT 2463.230 126.990 2464.410 128.170 ;
        RECT 2461.630 -26.910 2462.810 -25.730 ;
        RECT 2463.230 -26.910 2464.410 -25.730 ;
        RECT 2461.630 -28.510 2462.810 -27.330 ;
        RECT 2463.230 -28.510 2464.410 -27.330 ;
        RECT 2641.630 3547.010 2642.810 3548.190 ;
        RECT 2643.230 3547.010 2644.410 3548.190 ;
        RECT 2641.630 3545.410 2642.810 3546.590 ;
        RECT 2643.230 3545.410 2644.410 3546.590 ;
        RECT 2641.630 3368.590 2642.810 3369.770 ;
        RECT 2643.230 3368.590 2644.410 3369.770 ;
        RECT 2641.630 3366.990 2642.810 3368.170 ;
        RECT 2643.230 3366.990 2644.410 3368.170 ;
        RECT 2641.630 3188.590 2642.810 3189.770 ;
        RECT 2643.230 3188.590 2644.410 3189.770 ;
        RECT 2641.630 3186.990 2642.810 3188.170 ;
        RECT 2643.230 3186.990 2644.410 3188.170 ;
        RECT 2641.630 3008.590 2642.810 3009.770 ;
        RECT 2643.230 3008.590 2644.410 3009.770 ;
        RECT 2641.630 3006.990 2642.810 3008.170 ;
        RECT 2643.230 3006.990 2644.410 3008.170 ;
        RECT 2641.630 2828.590 2642.810 2829.770 ;
        RECT 2643.230 2828.590 2644.410 2829.770 ;
        RECT 2641.630 2826.990 2642.810 2828.170 ;
        RECT 2643.230 2826.990 2644.410 2828.170 ;
        RECT 2641.630 2648.590 2642.810 2649.770 ;
        RECT 2643.230 2648.590 2644.410 2649.770 ;
        RECT 2641.630 2646.990 2642.810 2648.170 ;
        RECT 2643.230 2646.990 2644.410 2648.170 ;
        RECT 2641.630 2468.590 2642.810 2469.770 ;
        RECT 2643.230 2468.590 2644.410 2469.770 ;
        RECT 2641.630 2466.990 2642.810 2468.170 ;
        RECT 2643.230 2466.990 2644.410 2468.170 ;
        RECT 2641.630 2288.590 2642.810 2289.770 ;
        RECT 2643.230 2288.590 2644.410 2289.770 ;
        RECT 2641.630 2286.990 2642.810 2288.170 ;
        RECT 2643.230 2286.990 2644.410 2288.170 ;
        RECT 2641.630 2108.590 2642.810 2109.770 ;
        RECT 2643.230 2108.590 2644.410 2109.770 ;
        RECT 2641.630 2106.990 2642.810 2108.170 ;
        RECT 2643.230 2106.990 2644.410 2108.170 ;
        RECT 2641.630 1928.590 2642.810 1929.770 ;
        RECT 2643.230 1928.590 2644.410 1929.770 ;
        RECT 2641.630 1926.990 2642.810 1928.170 ;
        RECT 2643.230 1926.990 2644.410 1928.170 ;
        RECT 2641.630 1748.590 2642.810 1749.770 ;
        RECT 2643.230 1748.590 2644.410 1749.770 ;
        RECT 2641.630 1746.990 2642.810 1748.170 ;
        RECT 2643.230 1746.990 2644.410 1748.170 ;
        RECT 2641.630 1568.590 2642.810 1569.770 ;
        RECT 2643.230 1568.590 2644.410 1569.770 ;
        RECT 2641.630 1566.990 2642.810 1568.170 ;
        RECT 2643.230 1566.990 2644.410 1568.170 ;
        RECT 2641.630 1388.590 2642.810 1389.770 ;
        RECT 2643.230 1388.590 2644.410 1389.770 ;
        RECT 2641.630 1386.990 2642.810 1388.170 ;
        RECT 2643.230 1386.990 2644.410 1388.170 ;
        RECT 2641.630 1208.590 2642.810 1209.770 ;
        RECT 2643.230 1208.590 2644.410 1209.770 ;
        RECT 2641.630 1206.990 2642.810 1208.170 ;
        RECT 2643.230 1206.990 2644.410 1208.170 ;
        RECT 2641.630 1028.590 2642.810 1029.770 ;
        RECT 2643.230 1028.590 2644.410 1029.770 ;
        RECT 2641.630 1026.990 2642.810 1028.170 ;
        RECT 2643.230 1026.990 2644.410 1028.170 ;
        RECT 2641.630 848.590 2642.810 849.770 ;
        RECT 2643.230 848.590 2644.410 849.770 ;
        RECT 2641.630 846.990 2642.810 848.170 ;
        RECT 2643.230 846.990 2644.410 848.170 ;
        RECT 2641.630 668.590 2642.810 669.770 ;
        RECT 2643.230 668.590 2644.410 669.770 ;
        RECT 2641.630 666.990 2642.810 668.170 ;
        RECT 2643.230 666.990 2644.410 668.170 ;
        RECT 2641.630 488.590 2642.810 489.770 ;
        RECT 2643.230 488.590 2644.410 489.770 ;
        RECT 2641.630 486.990 2642.810 488.170 ;
        RECT 2643.230 486.990 2644.410 488.170 ;
        RECT 2641.630 308.590 2642.810 309.770 ;
        RECT 2643.230 308.590 2644.410 309.770 ;
        RECT 2641.630 306.990 2642.810 308.170 ;
        RECT 2643.230 306.990 2644.410 308.170 ;
        RECT 2641.630 128.590 2642.810 129.770 ;
        RECT 2643.230 128.590 2644.410 129.770 ;
        RECT 2641.630 126.990 2642.810 128.170 ;
        RECT 2643.230 126.990 2644.410 128.170 ;
        RECT 2641.630 -26.910 2642.810 -25.730 ;
        RECT 2643.230 -26.910 2644.410 -25.730 ;
        RECT 2641.630 -28.510 2642.810 -27.330 ;
        RECT 2643.230 -28.510 2644.410 -27.330 ;
        RECT 2821.630 3547.010 2822.810 3548.190 ;
        RECT 2823.230 3547.010 2824.410 3548.190 ;
        RECT 2821.630 3545.410 2822.810 3546.590 ;
        RECT 2823.230 3545.410 2824.410 3546.590 ;
        RECT 2821.630 3368.590 2822.810 3369.770 ;
        RECT 2823.230 3368.590 2824.410 3369.770 ;
        RECT 2821.630 3366.990 2822.810 3368.170 ;
        RECT 2823.230 3366.990 2824.410 3368.170 ;
        RECT 2821.630 3188.590 2822.810 3189.770 ;
        RECT 2823.230 3188.590 2824.410 3189.770 ;
        RECT 2821.630 3186.990 2822.810 3188.170 ;
        RECT 2823.230 3186.990 2824.410 3188.170 ;
        RECT 2821.630 3008.590 2822.810 3009.770 ;
        RECT 2823.230 3008.590 2824.410 3009.770 ;
        RECT 2821.630 3006.990 2822.810 3008.170 ;
        RECT 2823.230 3006.990 2824.410 3008.170 ;
        RECT 2821.630 2828.590 2822.810 2829.770 ;
        RECT 2823.230 2828.590 2824.410 2829.770 ;
        RECT 2821.630 2826.990 2822.810 2828.170 ;
        RECT 2823.230 2826.990 2824.410 2828.170 ;
        RECT 2821.630 2648.590 2822.810 2649.770 ;
        RECT 2823.230 2648.590 2824.410 2649.770 ;
        RECT 2821.630 2646.990 2822.810 2648.170 ;
        RECT 2823.230 2646.990 2824.410 2648.170 ;
        RECT 2821.630 2468.590 2822.810 2469.770 ;
        RECT 2823.230 2468.590 2824.410 2469.770 ;
        RECT 2821.630 2466.990 2822.810 2468.170 ;
        RECT 2823.230 2466.990 2824.410 2468.170 ;
        RECT 2821.630 2288.590 2822.810 2289.770 ;
        RECT 2823.230 2288.590 2824.410 2289.770 ;
        RECT 2821.630 2286.990 2822.810 2288.170 ;
        RECT 2823.230 2286.990 2824.410 2288.170 ;
        RECT 2821.630 2108.590 2822.810 2109.770 ;
        RECT 2823.230 2108.590 2824.410 2109.770 ;
        RECT 2821.630 2106.990 2822.810 2108.170 ;
        RECT 2823.230 2106.990 2824.410 2108.170 ;
        RECT 2821.630 1928.590 2822.810 1929.770 ;
        RECT 2823.230 1928.590 2824.410 1929.770 ;
        RECT 2821.630 1926.990 2822.810 1928.170 ;
        RECT 2823.230 1926.990 2824.410 1928.170 ;
        RECT 2821.630 1748.590 2822.810 1749.770 ;
        RECT 2823.230 1748.590 2824.410 1749.770 ;
        RECT 2821.630 1746.990 2822.810 1748.170 ;
        RECT 2823.230 1746.990 2824.410 1748.170 ;
        RECT 2821.630 1568.590 2822.810 1569.770 ;
        RECT 2823.230 1568.590 2824.410 1569.770 ;
        RECT 2821.630 1566.990 2822.810 1568.170 ;
        RECT 2823.230 1566.990 2824.410 1568.170 ;
        RECT 2821.630 1388.590 2822.810 1389.770 ;
        RECT 2823.230 1388.590 2824.410 1389.770 ;
        RECT 2821.630 1386.990 2822.810 1388.170 ;
        RECT 2823.230 1386.990 2824.410 1388.170 ;
        RECT 2821.630 1208.590 2822.810 1209.770 ;
        RECT 2823.230 1208.590 2824.410 1209.770 ;
        RECT 2821.630 1206.990 2822.810 1208.170 ;
        RECT 2823.230 1206.990 2824.410 1208.170 ;
        RECT 2821.630 1028.590 2822.810 1029.770 ;
        RECT 2823.230 1028.590 2824.410 1029.770 ;
        RECT 2821.630 1026.990 2822.810 1028.170 ;
        RECT 2823.230 1026.990 2824.410 1028.170 ;
        RECT 2821.630 848.590 2822.810 849.770 ;
        RECT 2823.230 848.590 2824.410 849.770 ;
        RECT 2821.630 846.990 2822.810 848.170 ;
        RECT 2823.230 846.990 2824.410 848.170 ;
        RECT 2821.630 668.590 2822.810 669.770 ;
        RECT 2823.230 668.590 2824.410 669.770 ;
        RECT 2821.630 666.990 2822.810 668.170 ;
        RECT 2823.230 666.990 2824.410 668.170 ;
        RECT 2821.630 488.590 2822.810 489.770 ;
        RECT 2823.230 488.590 2824.410 489.770 ;
        RECT 2821.630 486.990 2822.810 488.170 ;
        RECT 2823.230 486.990 2824.410 488.170 ;
        RECT 2821.630 308.590 2822.810 309.770 ;
        RECT 2823.230 308.590 2824.410 309.770 ;
        RECT 2821.630 306.990 2822.810 308.170 ;
        RECT 2823.230 306.990 2824.410 308.170 ;
        RECT 2821.630 128.590 2822.810 129.770 ;
        RECT 2823.230 128.590 2824.410 129.770 ;
        RECT 2821.630 126.990 2822.810 128.170 ;
        RECT 2823.230 126.990 2824.410 128.170 ;
        RECT 2821.630 -26.910 2822.810 -25.730 ;
        RECT 2823.230 -26.910 2824.410 -25.730 ;
        RECT 2821.630 -28.510 2822.810 -27.330 ;
        RECT 2823.230 -28.510 2824.410 -27.330 ;
        RECT 2950.710 3547.010 2951.890 3548.190 ;
        RECT 2952.310 3547.010 2953.490 3548.190 ;
        RECT 2950.710 3545.410 2951.890 3546.590 ;
        RECT 2952.310 3545.410 2953.490 3546.590 ;
        RECT 2950.710 3368.590 2951.890 3369.770 ;
        RECT 2952.310 3368.590 2953.490 3369.770 ;
        RECT 2950.710 3366.990 2951.890 3368.170 ;
        RECT 2952.310 3366.990 2953.490 3368.170 ;
        RECT 2950.710 3188.590 2951.890 3189.770 ;
        RECT 2952.310 3188.590 2953.490 3189.770 ;
        RECT 2950.710 3186.990 2951.890 3188.170 ;
        RECT 2952.310 3186.990 2953.490 3188.170 ;
        RECT 2950.710 3008.590 2951.890 3009.770 ;
        RECT 2952.310 3008.590 2953.490 3009.770 ;
        RECT 2950.710 3006.990 2951.890 3008.170 ;
        RECT 2952.310 3006.990 2953.490 3008.170 ;
        RECT 2950.710 2828.590 2951.890 2829.770 ;
        RECT 2952.310 2828.590 2953.490 2829.770 ;
        RECT 2950.710 2826.990 2951.890 2828.170 ;
        RECT 2952.310 2826.990 2953.490 2828.170 ;
        RECT 2950.710 2648.590 2951.890 2649.770 ;
        RECT 2952.310 2648.590 2953.490 2649.770 ;
        RECT 2950.710 2646.990 2951.890 2648.170 ;
        RECT 2952.310 2646.990 2953.490 2648.170 ;
        RECT 2950.710 2468.590 2951.890 2469.770 ;
        RECT 2952.310 2468.590 2953.490 2469.770 ;
        RECT 2950.710 2466.990 2951.890 2468.170 ;
        RECT 2952.310 2466.990 2953.490 2468.170 ;
        RECT 2950.710 2288.590 2951.890 2289.770 ;
        RECT 2952.310 2288.590 2953.490 2289.770 ;
        RECT 2950.710 2286.990 2951.890 2288.170 ;
        RECT 2952.310 2286.990 2953.490 2288.170 ;
        RECT 2950.710 2108.590 2951.890 2109.770 ;
        RECT 2952.310 2108.590 2953.490 2109.770 ;
        RECT 2950.710 2106.990 2951.890 2108.170 ;
        RECT 2952.310 2106.990 2953.490 2108.170 ;
        RECT 2950.710 1928.590 2951.890 1929.770 ;
        RECT 2952.310 1928.590 2953.490 1929.770 ;
        RECT 2950.710 1926.990 2951.890 1928.170 ;
        RECT 2952.310 1926.990 2953.490 1928.170 ;
        RECT 2950.710 1748.590 2951.890 1749.770 ;
        RECT 2952.310 1748.590 2953.490 1749.770 ;
        RECT 2950.710 1746.990 2951.890 1748.170 ;
        RECT 2952.310 1746.990 2953.490 1748.170 ;
        RECT 2950.710 1568.590 2951.890 1569.770 ;
        RECT 2952.310 1568.590 2953.490 1569.770 ;
        RECT 2950.710 1566.990 2951.890 1568.170 ;
        RECT 2952.310 1566.990 2953.490 1568.170 ;
        RECT 2950.710 1388.590 2951.890 1389.770 ;
        RECT 2952.310 1388.590 2953.490 1389.770 ;
        RECT 2950.710 1386.990 2951.890 1388.170 ;
        RECT 2952.310 1386.990 2953.490 1388.170 ;
        RECT 2950.710 1208.590 2951.890 1209.770 ;
        RECT 2952.310 1208.590 2953.490 1209.770 ;
        RECT 2950.710 1206.990 2951.890 1208.170 ;
        RECT 2952.310 1206.990 2953.490 1208.170 ;
        RECT 2950.710 1028.590 2951.890 1029.770 ;
        RECT 2952.310 1028.590 2953.490 1029.770 ;
        RECT 2950.710 1026.990 2951.890 1028.170 ;
        RECT 2952.310 1026.990 2953.490 1028.170 ;
        RECT 2950.710 848.590 2951.890 849.770 ;
        RECT 2952.310 848.590 2953.490 849.770 ;
        RECT 2950.710 846.990 2951.890 848.170 ;
        RECT 2952.310 846.990 2953.490 848.170 ;
        RECT 2950.710 668.590 2951.890 669.770 ;
        RECT 2952.310 668.590 2953.490 669.770 ;
        RECT 2950.710 666.990 2951.890 668.170 ;
        RECT 2952.310 666.990 2953.490 668.170 ;
        RECT 2950.710 488.590 2951.890 489.770 ;
        RECT 2952.310 488.590 2953.490 489.770 ;
        RECT 2950.710 486.990 2951.890 488.170 ;
        RECT 2952.310 486.990 2953.490 488.170 ;
        RECT 2950.710 308.590 2951.890 309.770 ;
        RECT 2952.310 308.590 2953.490 309.770 ;
        RECT 2950.710 306.990 2951.890 308.170 ;
        RECT 2952.310 306.990 2953.490 308.170 ;
        RECT 2950.710 128.590 2951.890 129.770 ;
        RECT 2952.310 128.590 2953.490 129.770 ;
        RECT 2950.710 126.990 2951.890 128.170 ;
        RECT 2952.310 126.990 2953.490 128.170 ;
        RECT 2950.710 -26.910 2951.890 -25.730 ;
        RECT 2952.310 -26.910 2953.490 -25.730 ;
        RECT 2950.710 -28.510 2951.890 -27.330 ;
        RECT 2952.310 -28.510 2953.490 -27.330 ;
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
        RECT -43.630 3366.830 2963.250 3369.930 ;
        RECT -43.630 3186.830 2963.250 3189.930 ;
        RECT -43.630 3006.830 2963.250 3009.930 ;
        RECT -43.630 2826.830 2963.250 2829.930 ;
        RECT -43.630 2646.830 2963.250 2649.930 ;
        RECT -43.630 2466.830 2963.250 2469.930 ;
        RECT -43.630 2286.830 2963.250 2289.930 ;
        RECT -43.630 2106.830 2963.250 2109.930 ;
        RECT -43.630 1926.830 2963.250 1929.930 ;
        RECT -43.630 1746.830 2963.250 1749.930 ;
        RECT -43.630 1566.830 2963.250 1569.930 ;
        RECT -43.630 1386.830 2963.250 1389.930 ;
        RECT -43.630 1206.830 2963.250 1209.930 ;
        RECT -43.630 1026.830 2963.250 1029.930 ;
        RECT -43.630 846.830 2963.250 849.930 ;
        RECT -43.630 666.830 2963.250 669.930 ;
        RECT -43.630 486.830 2963.250 489.930 ;
        RECT -43.630 306.830 2963.250 309.930 ;
        RECT -43.630 126.830 2963.250 129.930 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
        RECT 166.470 -38.270 169.570 3557.950 ;
        RECT 346.470 -38.270 349.570 3557.950 ;
        RECT 526.470 810.000 529.570 3557.950 ;
        RECT 706.470 810.000 709.570 3557.950 ;
        RECT 526.470 -38.270 529.570 490.000 ;
        RECT 706.470 -38.270 709.570 490.000 ;
        RECT 886.470 -38.270 889.570 3557.950 ;
        RECT 1066.470 -38.270 1069.570 3557.950 ;
        RECT 1246.470 -38.270 1249.570 3557.950 ;
        RECT 1426.470 -38.270 1429.570 3557.950 ;
        RECT 1606.470 -38.270 1609.570 3557.950 ;
        RECT 1786.470 -38.270 1789.570 3557.950 ;
        RECT 1966.470 -38.270 1969.570 3557.950 ;
        RECT 2146.470 -38.270 2149.570 3557.950 ;
        RECT 2326.470 -38.270 2329.570 3557.950 ;
        RECT 2506.470 -38.270 2509.570 3557.950 ;
        RECT 2686.470 -38.270 2689.570 3557.950 ;
        RECT 2866.470 -38.270 2869.570 3557.950 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
      LAYER via4 ;
        RECT -43.470 3556.610 -42.290 3557.790 ;
        RECT -41.870 3556.610 -40.690 3557.790 ;
        RECT -43.470 3555.010 -42.290 3556.190 ;
        RECT -41.870 3555.010 -40.690 3556.190 ;
        RECT -43.470 3413.590 -42.290 3414.770 ;
        RECT -41.870 3413.590 -40.690 3414.770 ;
        RECT -43.470 3411.990 -42.290 3413.170 ;
        RECT -41.870 3411.990 -40.690 3413.170 ;
        RECT -43.470 3233.590 -42.290 3234.770 ;
        RECT -41.870 3233.590 -40.690 3234.770 ;
        RECT -43.470 3231.990 -42.290 3233.170 ;
        RECT -41.870 3231.990 -40.690 3233.170 ;
        RECT -43.470 3053.590 -42.290 3054.770 ;
        RECT -41.870 3053.590 -40.690 3054.770 ;
        RECT -43.470 3051.990 -42.290 3053.170 ;
        RECT -41.870 3051.990 -40.690 3053.170 ;
        RECT -43.470 2873.590 -42.290 2874.770 ;
        RECT -41.870 2873.590 -40.690 2874.770 ;
        RECT -43.470 2871.990 -42.290 2873.170 ;
        RECT -41.870 2871.990 -40.690 2873.170 ;
        RECT -43.470 2693.590 -42.290 2694.770 ;
        RECT -41.870 2693.590 -40.690 2694.770 ;
        RECT -43.470 2691.990 -42.290 2693.170 ;
        RECT -41.870 2691.990 -40.690 2693.170 ;
        RECT -43.470 2513.590 -42.290 2514.770 ;
        RECT -41.870 2513.590 -40.690 2514.770 ;
        RECT -43.470 2511.990 -42.290 2513.170 ;
        RECT -41.870 2511.990 -40.690 2513.170 ;
        RECT -43.470 2333.590 -42.290 2334.770 ;
        RECT -41.870 2333.590 -40.690 2334.770 ;
        RECT -43.470 2331.990 -42.290 2333.170 ;
        RECT -41.870 2331.990 -40.690 2333.170 ;
        RECT -43.470 2153.590 -42.290 2154.770 ;
        RECT -41.870 2153.590 -40.690 2154.770 ;
        RECT -43.470 2151.990 -42.290 2153.170 ;
        RECT -41.870 2151.990 -40.690 2153.170 ;
        RECT -43.470 1973.590 -42.290 1974.770 ;
        RECT -41.870 1973.590 -40.690 1974.770 ;
        RECT -43.470 1971.990 -42.290 1973.170 ;
        RECT -41.870 1971.990 -40.690 1973.170 ;
        RECT -43.470 1793.590 -42.290 1794.770 ;
        RECT -41.870 1793.590 -40.690 1794.770 ;
        RECT -43.470 1791.990 -42.290 1793.170 ;
        RECT -41.870 1791.990 -40.690 1793.170 ;
        RECT -43.470 1613.590 -42.290 1614.770 ;
        RECT -41.870 1613.590 -40.690 1614.770 ;
        RECT -43.470 1611.990 -42.290 1613.170 ;
        RECT -41.870 1611.990 -40.690 1613.170 ;
        RECT -43.470 1433.590 -42.290 1434.770 ;
        RECT -41.870 1433.590 -40.690 1434.770 ;
        RECT -43.470 1431.990 -42.290 1433.170 ;
        RECT -41.870 1431.990 -40.690 1433.170 ;
        RECT -43.470 1253.590 -42.290 1254.770 ;
        RECT -41.870 1253.590 -40.690 1254.770 ;
        RECT -43.470 1251.990 -42.290 1253.170 ;
        RECT -41.870 1251.990 -40.690 1253.170 ;
        RECT -43.470 1073.590 -42.290 1074.770 ;
        RECT -41.870 1073.590 -40.690 1074.770 ;
        RECT -43.470 1071.990 -42.290 1073.170 ;
        RECT -41.870 1071.990 -40.690 1073.170 ;
        RECT -43.470 893.590 -42.290 894.770 ;
        RECT -41.870 893.590 -40.690 894.770 ;
        RECT -43.470 891.990 -42.290 893.170 ;
        RECT -41.870 891.990 -40.690 893.170 ;
        RECT -43.470 713.590 -42.290 714.770 ;
        RECT -41.870 713.590 -40.690 714.770 ;
        RECT -43.470 711.990 -42.290 713.170 ;
        RECT -41.870 711.990 -40.690 713.170 ;
        RECT -43.470 533.590 -42.290 534.770 ;
        RECT -41.870 533.590 -40.690 534.770 ;
        RECT -43.470 531.990 -42.290 533.170 ;
        RECT -41.870 531.990 -40.690 533.170 ;
        RECT -43.470 353.590 -42.290 354.770 ;
        RECT -41.870 353.590 -40.690 354.770 ;
        RECT -43.470 351.990 -42.290 353.170 ;
        RECT -41.870 351.990 -40.690 353.170 ;
        RECT -43.470 173.590 -42.290 174.770 ;
        RECT -41.870 173.590 -40.690 174.770 ;
        RECT -43.470 171.990 -42.290 173.170 ;
        RECT -41.870 171.990 -40.690 173.170 ;
        RECT -43.470 -36.510 -42.290 -35.330 ;
        RECT -41.870 -36.510 -40.690 -35.330 ;
        RECT -43.470 -38.110 -42.290 -36.930 ;
        RECT -41.870 -38.110 -40.690 -36.930 ;
        RECT 166.630 3556.610 167.810 3557.790 ;
        RECT 168.230 3556.610 169.410 3557.790 ;
        RECT 166.630 3555.010 167.810 3556.190 ;
        RECT 168.230 3555.010 169.410 3556.190 ;
        RECT 166.630 3413.590 167.810 3414.770 ;
        RECT 168.230 3413.590 169.410 3414.770 ;
        RECT 166.630 3411.990 167.810 3413.170 ;
        RECT 168.230 3411.990 169.410 3413.170 ;
        RECT 166.630 3233.590 167.810 3234.770 ;
        RECT 168.230 3233.590 169.410 3234.770 ;
        RECT 166.630 3231.990 167.810 3233.170 ;
        RECT 168.230 3231.990 169.410 3233.170 ;
        RECT 166.630 3053.590 167.810 3054.770 ;
        RECT 168.230 3053.590 169.410 3054.770 ;
        RECT 166.630 3051.990 167.810 3053.170 ;
        RECT 168.230 3051.990 169.410 3053.170 ;
        RECT 166.630 2873.590 167.810 2874.770 ;
        RECT 168.230 2873.590 169.410 2874.770 ;
        RECT 166.630 2871.990 167.810 2873.170 ;
        RECT 168.230 2871.990 169.410 2873.170 ;
        RECT 166.630 2693.590 167.810 2694.770 ;
        RECT 168.230 2693.590 169.410 2694.770 ;
        RECT 166.630 2691.990 167.810 2693.170 ;
        RECT 168.230 2691.990 169.410 2693.170 ;
        RECT 166.630 2513.590 167.810 2514.770 ;
        RECT 168.230 2513.590 169.410 2514.770 ;
        RECT 166.630 2511.990 167.810 2513.170 ;
        RECT 168.230 2511.990 169.410 2513.170 ;
        RECT 166.630 2333.590 167.810 2334.770 ;
        RECT 168.230 2333.590 169.410 2334.770 ;
        RECT 166.630 2331.990 167.810 2333.170 ;
        RECT 168.230 2331.990 169.410 2333.170 ;
        RECT 166.630 2153.590 167.810 2154.770 ;
        RECT 168.230 2153.590 169.410 2154.770 ;
        RECT 166.630 2151.990 167.810 2153.170 ;
        RECT 168.230 2151.990 169.410 2153.170 ;
        RECT 166.630 1973.590 167.810 1974.770 ;
        RECT 168.230 1973.590 169.410 1974.770 ;
        RECT 166.630 1971.990 167.810 1973.170 ;
        RECT 168.230 1971.990 169.410 1973.170 ;
        RECT 166.630 1793.590 167.810 1794.770 ;
        RECT 168.230 1793.590 169.410 1794.770 ;
        RECT 166.630 1791.990 167.810 1793.170 ;
        RECT 168.230 1791.990 169.410 1793.170 ;
        RECT 166.630 1613.590 167.810 1614.770 ;
        RECT 168.230 1613.590 169.410 1614.770 ;
        RECT 166.630 1611.990 167.810 1613.170 ;
        RECT 168.230 1611.990 169.410 1613.170 ;
        RECT 166.630 1433.590 167.810 1434.770 ;
        RECT 168.230 1433.590 169.410 1434.770 ;
        RECT 166.630 1431.990 167.810 1433.170 ;
        RECT 168.230 1431.990 169.410 1433.170 ;
        RECT 166.630 1253.590 167.810 1254.770 ;
        RECT 168.230 1253.590 169.410 1254.770 ;
        RECT 166.630 1251.990 167.810 1253.170 ;
        RECT 168.230 1251.990 169.410 1253.170 ;
        RECT 166.630 1073.590 167.810 1074.770 ;
        RECT 168.230 1073.590 169.410 1074.770 ;
        RECT 166.630 1071.990 167.810 1073.170 ;
        RECT 168.230 1071.990 169.410 1073.170 ;
        RECT 166.630 893.590 167.810 894.770 ;
        RECT 168.230 893.590 169.410 894.770 ;
        RECT 166.630 891.990 167.810 893.170 ;
        RECT 168.230 891.990 169.410 893.170 ;
        RECT 166.630 713.590 167.810 714.770 ;
        RECT 168.230 713.590 169.410 714.770 ;
        RECT 166.630 711.990 167.810 713.170 ;
        RECT 168.230 711.990 169.410 713.170 ;
        RECT 166.630 533.590 167.810 534.770 ;
        RECT 168.230 533.590 169.410 534.770 ;
        RECT 166.630 531.990 167.810 533.170 ;
        RECT 168.230 531.990 169.410 533.170 ;
        RECT 166.630 353.590 167.810 354.770 ;
        RECT 168.230 353.590 169.410 354.770 ;
        RECT 166.630 351.990 167.810 353.170 ;
        RECT 168.230 351.990 169.410 353.170 ;
        RECT 166.630 173.590 167.810 174.770 ;
        RECT 168.230 173.590 169.410 174.770 ;
        RECT 166.630 171.990 167.810 173.170 ;
        RECT 168.230 171.990 169.410 173.170 ;
        RECT 166.630 -36.510 167.810 -35.330 ;
        RECT 168.230 -36.510 169.410 -35.330 ;
        RECT 166.630 -38.110 167.810 -36.930 ;
        RECT 168.230 -38.110 169.410 -36.930 ;
        RECT 346.630 3556.610 347.810 3557.790 ;
        RECT 348.230 3556.610 349.410 3557.790 ;
        RECT 346.630 3555.010 347.810 3556.190 ;
        RECT 348.230 3555.010 349.410 3556.190 ;
        RECT 346.630 3413.590 347.810 3414.770 ;
        RECT 348.230 3413.590 349.410 3414.770 ;
        RECT 346.630 3411.990 347.810 3413.170 ;
        RECT 348.230 3411.990 349.410 3413.170 ;
        RECT 346.630 3233.590 347.810 3234.770 ;
        RECT 348.230 3233.590 349.410 3234.770 ;
        RECT 346.630 3231.990 347.810 3233.170 ;
        RECT 348.230 3231.990 349.410 3233.170 ;
        RECT 346.630 3053.590 347.810 3054.770 ;
        RECT 348.230 3053.590 349.410 3054.770 ;
        RECT 346.630 3051.990 347.810 3053.170 ;
        RECT 348.230 3051.990 349.410 3053.170 ;
        RECT 346.630 2873.590 347.810 2874.770 ;
        RECT 348.230 2873.590 349.410 2874.770 ;
        RECT 346.630 2871.990 347.810 2873.170 ;
        RECT 348.230 2871.990 349.410 2873.170 ;
        RECT 346.630 2693.590 347.810 2694.770 ;
        RECT 348.230 2693.590 349.410 2694.770 ;
        RECT 346.630 2691.990 347.810 2693.170 ;
        RECT 348.230 2691.990 349.410 2693.170 ;
        RECT 346.630 2513.590 347.810 2514.770 ;
        RECT 348.230 2513.590 349.410 2514.770 ;
        RECT 346.630 2511.990 347.810 2513.170 ;
        RECT 348.230 2511.990 349.410 2513.170 ;
        RECT 346.630 2333.590 347.810 2334.770 ;
        RECT 348.230 2333.590 349.410 2334.770 ;
        RECT 346.630 2331.990 347.810 2333.170 ;
        RECT 348.230 2331.990 349.410 2333.170 ;
        RECT 346.630 2153.590 347.810 2154.770 ;
        RECT 348.230 2153.590 349.410 2154.770 ;
        RECT 346.630 2151.990 347.810 2153.170 ;
        RECT 348.230 2151.990 349.410 2153.170 ;
        RECT 346.630 1973.590 347.810 1974.770 ;
        RECT 348.230 1973.590 349.410 1974.770 ;
        RECT 346.630 1971.990 347.810 1973.170 ;
        RECT 348.230 1971.990 349.410 1973.170 ;
        RECT 346.630 1793.590 347.810 1794.770 ;
        RECT 348.230 1793.590 349.410 1794.770 ;
        RECT 346.630 1791.990 347.810 1793.170 ;
        RECT 348.230 1791.990 349.410 1793.170 ;
        RECT 346.630 1613.590 347.810 1614.770 ;
        RECT 348.230 1613.590 349.410 1614.770 ;
        RECT 346.630 1611.990 347.810 1613.170 ;
        RECT 348.230 1611.990 349.410 1613.170 ;
        RECT 346.630 1433.590 347.810 1434.770 ;
        RECT 348.230 1433.590 349.410 1434.770 ;
        RECT 346.630 1431.990 347.810 1433.170 ;
        RECT 348.230 1431.990 349.410 1433.170 ;
        RECT 346.630 1253.590 347.810 1254.770 ;
        RECT 348.230 1253.590 349.410 1254.770 ;
        RECT 346.630 1251.990 347.810 1253.170 ;
        RECT 348.230 1251.990 349.410 1253.170 ;
        RECT 346.630 1073.590 347.810 1074.770 ;
        RECT 348.230 1073.590 349.410 1074.770 ;
        RECT 346.630 1071.990 347.810 1073.170 ;
        RECT 348.230 1071.990 349.410 1073.170 ;
        RECT 346.630 893.590 347.810 894.770 ;
        RECT 348.230 893.590 349.410 894.770 ;
        RECT 346.630 891.990 347.810 893.170 ;
        RECT 348.230 891.990 349.410 893.170 ;
        RECT 526.630 3556.610 527.810 3557.790 ;
        RECT 528.230 3556.610 529.410 3557.790 ;
        RECT 526.630 3555.010 527.810 3556.190 ;
        RECT 528.230 3555.010 529.410 3556.190 ;
        RECT 526.630 3413.590 527.810 3414.770 ;
        RECT 528.230 3413.590 529.410 3414.770 ;
        RECT 526.630 3411.990 527.810 3413.170 ;
        RECT 528.230 3411.990 529.410 3413.170 ;
        RECT 526.630 3233.590 527.810 3234.770 ;
        RECT 528.230 3233.590 529.410 3234.770 ;
        RECT 526.630 3231.990 527.810 3233.170 ;
        RECT 528.230 3231.990 529.410 3233.170 ;
        RECT 526.630 3053.590 527.810 3054.770 ;
        RECT 528.230 3053.590 529.410 3054.770 ;
        RECT 526.630 3051.990 527.810 3053.170 ;
        RECT 528.230 3051.990 529.410 3053.170 ;
        RECT 526.630 2873.590 527.810 2874.770 ;
        RECT 528.230 2873.590 529.410 2874.770 ;
        RECT 526.630 2871.990 527.810 2873.170 ;
        RECT 528.230 2871.990 529.410 2873.170 ;
        RECT 526.630 2693.590 527.810 2694.770 ;
        RECT 528.230 2693.590 529.410 2694.770 ;
        RECT 526.630 2691.990 527.810 2693.170 ;
        RECT 528.230 2691.990 529.410 2693.170 ;
        RECT 526.630 2513.590 527.810 2514.770 ;
        RECT 528.230 2513.590 529.410 2514.770 ;
        RECT 526.630 2511.990 527.810 2513.170 ;
        RECT 528.230 2511.990 529.410 2513.170 ;
        RECT 526.630 2333.590 527.810 2334.770 ;
        RECT 528.230 2333.590 529.410 2334.770 ;
        RECT 526.630 2331.990 527.810 2333.170 ;
        RECT 528.230 2331.990 529.410 2333.170 ;
        RECT 526.630 2153.590 527.810 2154.770 ;
        RECT 528.230 2153.590 529.410 2154.770 ;
        RECT 526.630 2151.990 527.810 2153.170 ;
        RECT 528.230 2151.990 529.410 2153.170 ;
        RECT 526.630 1973.590 527.810 1974.770 ;
        RECT 528.230 1973.590 529.410 1974.770 ;
        RECT 526.630 1971.990 527.810 1973.170 ;
        RECT 528.230 1971.990 529.410 1973.170 ;
        RECT 526.630 1793.590 527.810 1794.770 ;
        RECT 528.230 1793.590 529.410 1794.770 ;
        RECT 526.630 1791.990 527.810 1793.170 ;
        RECT 528.230 1791.990 529.410 1793.170 ;
        RECT 526.630 1613.590 527.810 1614.770 ;
        RECT 528.230 1613.590 529.410 1614.770 ;
        RECT 526.630 1611.990 527.810 1613.170 ;
        RECT 528.230 1611.990 529.410 1613.170 ;
        RECT 526.630 1433.590 527.810 1434.770 ;
        RECT 528.230 1433.590 529.410 1434.770 ;
        RECT 526.630 1431.990 527.810 1433.170 ;
        RECT 528.230 1431.990 529.410 1433.170 ;
        RECT 526.630 1253.590 527.810 1254.770 ;
        RECT 528.230 1253.590 529.410 1254.770 ;
        RECT 526.630 1251.990 527.810 1253.170 ;
        RECT 528.230 1251.990 529.410 1253.170 ;
        RECT 526.630 1073.590 527.810 1074.770 ;
        RECT 528.230 1073.590 529.410 1074.770 ;
        RECT 526.630 1071.990 527.810 1073.170 ;
        RECT 528.230 1071.990 529.410 1073.170 ;
        RECT 526.630 893.590 527.810 894.770 ;
        RECT 528.230 893.590 529.410 894.770 ;
        RECT 526.630 891.990 527.810 893.170 ;
        RECT 528.230 891.990 529.410 893.170 ;
        RECT 706.630 3556.610 707.810 3557.790 ;
        RECT 708.230 3556.610 709.410 3557.790 ;
        RECT 706.630 3555.010 707.810 3556.190 ;
        RECT 708.230 3555.010 709.410 3556.190 ;
        RECT 706.630 3413.590 707.810 3414.770 ;
        RECT 708.230 3413.590 709.410 3414.770 ;
        RECT 706.630 3411.990 707.810 3413.170 ;
        RECT 708.230 3411.990 709.410 3413.170 ;
        RECT 706.630 3233.590 707.810 3234.770 ;
        RECT 708.230 3233.590 709.410 3234.770 ;
        RECT 706.630 3231.990 707.810 3233.170 ;
        RECT 708.230 3231.990 709.410 3233.170 ;
        RECT 706.630 3053.590 707.810 3054.770 ;
        RECT 708.230 3053.590 709.410 3054.770 ;
        RECT 706.630 3051.990 707.810 3053.170 ;
        RECT 708.230 3051.990 709.410 3053.170 ;
        RECT 706.630 2873.590 707.810 2874.770 ;
        RECT 708.230 2873.590 709.410 2874.770 ;
        RECT 706.630 2871.990 707.810 2873.170 ;
        RECT 708.230 2871.990 709.410 2873.170 ;
        RECT 706.630 2693.590 707.810 2694.770 ;
        RECT 708.230 2693.590 709.410 2694.770 ;
        RECT 706.630 2691.990 707.810 2693.170 ;
        RECT 708.230 2691.990 709.410 2693.170 ;
        RECT 706.630 2513.590 707.810 2514.770 ;
        RECT 708.230 2513.590 709.410 2514.770 ;
        RECT 706.630 2511.990 707.810 2513.170 ;
        RECT 708.230 2511.990 709.410 2513.170 ;
        RECT 706.630 2333.590 707.810 2334.770 ;
        RECT 708.230 2333.590 709.410 2334.770 ;
        RECT 706.630 2331.990 707.810 2333.170 ;
        RECT 708.230 2331.990 709.410 2333.170 ;
        RECT 706.630 2153.590 707.810 2154.770 ;
        RECT 708.230 2153.590 709.410 2154.770 ;
        RECT 706.630 2151.990 707.810 2153.170 ;
        RECT 708.230 2151.990 709.410 2153.170 ;
        RECT 706.630 1973.590 707.810 1974.770 ;
        RECT 708.230 1973.590 709.410 1974.770 ;
        RECT 706.630 1971.990 707.810 1973.170 ;
        RECT 708.230 1971.990 709.410 1973.170 ;
        RECT 706.630 1793.590 707.810 1794.770 ;
        RECT 708.230 1793.590 709.410 1794.770 ;
        RECT 706.630 1791.990 707.810 1793.170 ;
        RECT 708.230 1791.990 709.410 1793.170 ;
        RECT 706.630 1613.590 707.810 1614.770 ;
        RECT 708.230 1613.590 709.410 1614.770 ;
        RECT 706.630 1611.990 707.810 1613.170 ;
        RECT 708.230 1611.990 709.410 1613.170 ;
        RECT 706.630 1433.590 707.810 1434.770 ;
        RECT 708.230 1433.590 709.410 1434.770 ;
        RECT 706.630 1431.990 707.810 1433.170 ;
        RECT 708.230 1431.990 709.410 1433.170 ;
        RECT 706.630 1253.590 707.810 1254.770 ;
        RECT 708.230 1253.590 709.410 1254.770 ;
        RECT 706.630 1251.990 707.810 1253.170 ;
        RECT 708.230 1251.990 709.410 1253.170 ;
        RECT 706.630 1073.590 707.810 1074.770 ;
        RECT 708.230 1073.590 709.410 1074.770 ;
        RECT 706.630 1071.990 707.810 1073.170 ;
        RECT 708.230 1071.990 709.410 1073.170 ;
        RECT 706.630 893.590 707.810 894.770 ;
        RECT 708.230 893.590 709.410 894.770 ;
        RECT 706.630 891.990 707.810 893.170 ;
        RECT 708.230 891.990 709.410 893.170 ;
        RECT 886.630 3556.610 887.810 3557.790 ;
        RECT 888.230 3556.610 889.410 3557.790 ;
        RECT 886.630 3555.010 887.810 3556.190 ;
        RECT 888.230 3555.010 889.410 3556.190 ;
        RECT 886.630 3413.590 887.810 3414.770 ;
        RECT 888.230 3413.590 889.410 3414.770 ;
        RECT 886.630 3411.990 887.810 3413.170 ;
        RECT 888.230 3411.990 889.410 3413.170 ;
        RECT 886.630 3233.590 887.810 3234.770 ;
        RECT 888.230 3233.590 889.410 3234.770 ;
        RECT 886.630 3231.990 887.810 3233.170 ;
        RECT 888.230 3231.990 889.410 3233.170 ;
        RECT 886.630 3053.590 887.810 3054.770 ;
        RECT 888.230 3053.590 889.410 3054.770 ;
        RECT 886.630 3051.990 887.810 3053.170 ;
        RECT 888.230 3051.990 889.410 3053.170 ;
        RECT 886.630 2873.590 887.810 2874.770 ;
        RECT 888.230 2873.590 889.410 2874.770 ;
        RECT 886.630 2871.990 887.810 2873.170 ;
        RECT 888.230 2871.990 889.410 2873.170 ;
        RECT 886.630 2693.590 887.810 2694.770 ;
        RECT 888.230 2693.590 889.410 2694.770 ;
        RECT 886.630 2691.990 887.810 2693.170 ;
        RECT 888.230 2691.990 889.410 2693.170 ;
        RECT 886.630 2513.590 887.810 2514.770 ;
        RECT 888.230 2513.590 889.410 2514.770 ;
        RECT 886.630 2511.990 887.810 2513.170 ;
        RECT 888.230 2511.990 889.410 2513.170 ;
        RECT 886.630 2333.590 887.810 2334.770 ;
        RECT 888.230 2333.590 889.410 2334.770 ;
        RECT 886.630 2331.990 887.810 2333.170 ;
        RECT 888.230 2331.990 889.410 2333.170 ;
        RECT 886.630 2153.590 887.810 2154.770 ;
        RECT 888.230 2153.590 889.410 2154.770 ;
        RECT 886.630 2151.990 887.810 2153.170 ;
        RECT 888.230 2151.990 889.410 2153.170 ;
        RECT 886.630 1973.590 887.810 1974.770 ;
        RECT 888.230 1973.590 889.410 1974.770 ;
        RECT 886.630 1971.990 887.810 1973.170 ;
        RECT 888.230 1971.990 889.410 1973.170 ;
        RECT 886.630 1793.590 887.810 1794.770 ;
        RECT 888.230 1793.590 889.410 1794.770 ;
        RECT 886.630 1791.990 887.810 1793.170 ;
        RECT 888.230 1791.990 889.410 1793.170 ;
        RECT 886.630 1613.590 887.810 1614.770 ;
        RECT 888.230 1613.590 889.410 1614.770 ;
        RECT 886.630 1611.990 887.810 1613.170 ;
        RECT 888.230 1611.990 889.410 1613.170 ;
        RECT 886.630 1433.590 887.810 1434.770 ;
        RECT 888.230 1433.590 889.410 1434.770 ;
        RECT 886.630 1431.990 887.810 1433.170 ;
        RECT 888.230 1431.990 889.410 1433.170 ;
        RECT 886.630 1253.590 887.810 1254.770 ;
        RECT 888.230 1253.590 889.410 1254.770 ;
        RECT 886.630 1251.990 887.810 1253.170 ;
        RECT 888.230 1251.990 889.410 1253.170 ;
        RECT 886.630 1073.590 887.810 1074.770 ;
        RECT 888.230 1073.590 889.410 1074.770 ;
        RECT 886.630 1071.990 887.810 1073.170 ;
        RECT 888.230 1071.990 889.410 1073.170 ;
        RECT 886.630 893.590 887.810 894.770 ;
        RECT 888.230 893.590 889.410 894.770 ;
        RECT 886.630 891.990 887.810 893.170 ;
        RECT 888.230 891.990 889.410 893.170 ;
        RECT 346.630 713.590 347.810 714.770 ;
        RECT 348.230 713.590 349.410 714.770 ;
        RECT 346.630 711.990 347.810 713.170 ;
        RECT 348.230 711.990 349.410 713.170 ;
        RECT 346.630 533.590 347.810 534.770 ;
        RECT 348.230 533.590 349.410 534.770 ;
        RECT 346.630 531.990 347.810 533.170 ;
        RECT 348.230 531.990 349.410 533.170 ;
        RECT 886.630 713.590 887.810 714.770 ;
        RECT 888.230 713.590 889.410 714.770 ;
        RECT 886.630 711.990 887.810 713.170 ;
        RECT 888.230 711.990 889.410 713.170 ;
        RECT 886.630 533.590 887.810 534.770 ;
        RECT 888.230 533.590 889.410 534.770 ;
        RECT 886.630 531.990 887.810 533.170 ;
        RECT 888.230 531.990 889.410 533.170 ;
        RECT 346.630 353.590 347.810 354.770 ;
        RECT 348.230 353.590 349.410 354.770 ;
        RECT 346.630 351.990 347.810 353.170 ;
        RECT 348.230 351.990 349.410 353.170 ;
        RECT 346.630 173.590 347.810 174.770 ;
        RECT 348.230 173.590 349.410 174.770 ;
        RECT 346.630 171.990 347.810 173.170 ;
        RECT 348.230 171.990 349.410 173.170 ;
        RECT 346.630 -36.510 347.810 -35.330 ;
        RECT 348.230 -36.510 349.410 -35.330 ;
        RECT 346.630 -38.110 347.810 -36.930 ;
        RECT 348.230 -38.110 349.410 -36.930 ;
        RECT 526.630 353.590 527.810 354.770 ;
        RECT 528.230 353.590 529.410 354.770 ;
        RECT 526.630 351.990 527.810 353.170 ;
        RECT 528.230 351.990 529.410 353.170 ;
        RECT 526.630 173.590 527.810 174.770 ;
        RECT 528.230 173.590 529.410 174.770 ;
        RECT 526.630 171.990 527.810 173.170 ;
        RECT 528.230 171.990 529.410 173.170 ;
        RECT 526.630 -36.510 527.810 -35.330 ;
        RECT 528.230 -36.510 529.410 -35.330 ;
        RECT 526.630 -38.110 527.810 -36.930 ;
        RECT 528.230 -38.110 529.410 -36.930 ;
        RECT 706.630 353.590 707.810 354.770 ;
        RECT 708.230 353.590 709.410 354.770 ;
        RECT 706.630 351.990 707.810 353.170 ;
        RECT 708.230 351.990 709.410 353.170 ;
        RECT 706.630 173.590 707.810 174.770 ;
        RECT 708.230 173.590 709.410 174.770 ;
        RECT 706.630 171.990 707.810 173.170 ;
        RECT 708.230 171.990 709.410 173.170 ;
        RECT 706.630 -36.510 707.810 -35.330 ;
        RECT 708.230 -36.510 709.410 -35.330 ;
        RECT 706.630 -38.110 707.810 -36.930 ;
        RECT 708.230 -38.110 709.410 -36.930 ;
        RECT 886.630 353.590 887.810 354.770 ;
        RECT 888.230 353.590 889.410 354.770 ;
        RECT 886.630 351.990 887.810 353.170 ;
        RECT 888.230 351.990 889.410 353.170 ;
        RECT 886.630 173.590 887.810 174.770 ;
        RECT 888.230 173.590 889.410 174.770 ;
        RECT 886.630 171.990 887.810 173.170 ;
        RECT 888.230 171.990 889.410 173.170 ;
        RECT 886.630 -36.510 887.810 -35.330 ;
        RECT 888.230 -36.510 889.410 -35.330 ;
        RECT 886.630 -38.110 887.810 -36.930 ;
        RECT 888.230 -38.110 889.410 -36.930 ;
        RECT 1066.630 3556.610 1067.810 3557.790 ;
        RECT 1068.230 3556.610 1069.410 3557.790 ;
        RECT 1066.630 3555.010 1067.810 3556.190 ;
        RECT 1068.230 3555.010 1069.410 3556.190 ;
        RECT 1066.630 3413.590 1067.810 3414.770 ;
        RECT 1068.230 3413.590 1069.410 3414.770 ;
        RECT 1066.630 3411.990 1067.810 3413.170 ;
        RECT 1068.230 3411.990 1069.410 3413.170 ;
        RECT 1066.630 3233.590 1067.810 3234.770 ;
        RECT 1068.230 3233.590 1069.410 3234.770 ;
        RECT 1066.630 3231.990 1067.810 3233.170 ;
        RECT 1068.230 3231.990 1069.410 3233.170 ;
        RECT 1066.630 3053.590 1067.810 3054.770 ;
        RECT 1068.230 3053.590 1069.410 3054.770 ;
        RECT 1066.630 3051.990 1067.810 3053.170 ;
        RECT 1068.230 3051.990 1069.410 3053.170 ;
        RECT 1066.630 2873.590 1067.810 2874.770 ;
        RECT 1068.230 2873.590 1069.410 2874.770 ;
        RECT 1066.630 2871.990 1067.810 2873.170 ;
        RECT 1068.230 2871.990 1069.410 2873.170 ;
        RECT 1066.630 2693.590 1067.810 2694.770 ;
        RECT 1068.230 2693.590 1069.410 2694.770 ;
        RECT 1066.630 2691.990 1067.810 2693.170 ;
        RECT 1068.230 2691.990 1069.410 2693.170 ;
        RECT 1066.630 2513.590 1067.810 2514.770 ;
        RECT 1068.230 2513.590 1069.410 2514.770 ;
        RECT 1066.630 2511.990 1067.810 2513.170 ;
        RECT 1068.230 2511.990 1069.410 2513.170 ;
        RECT 1066.630 2333.590 1067.810 2334.770 ;
        RECT 1068.230 2333.590 1069.410 2334.770 ;
        RECT 1066.630 2331.990 1067.810 2333.170 ;
        RECT 1068.230 2331.990 1069.410 2333.170 ;
        RECT 1066.630 2153.590 1067.810 2154.770 ;
        RECT 1068.230 2153.590 1069.410 2154.770 ;
        RECT 1066.630 2151.990 1067.810 2153.170 ;
        RECT 1068.230 2151.990 1069.410 2153.170 ;
        RECT 1066.630 1973.590 1067.810 1974.770 ;
        RECT 1068.230 1973.590 1069.410 1974.770 ;
        RECT 1066.630 1971.990 1067.810 1973.170 ;
        RECT 1068.230 1971.990 1069.410 1973.170 ;
        RECT 1066.630 1793.590 1067.810 1794.770 ;
        RECT 1068.230 1793.590 1069.410 1794.770 ;
        RECT 1066.630 1791.990 1067.810 1793.170 ;
        RECT 1068.230 1791.990 1069.410 1793.170 ;
        RECT 1066.630 1613.590 1067.810 1614.770 ;
        RECT 1068.230 1613.590 1069.410 1614.770 ;
        RECT 1066.630 1611.990 1067.810 1613.170 ;
        RECT 1068.230 1611.990 1069.410 1613.170 ;
        RECT 1066.630 1433.590 1067.810 1434.770 ;
        RECT 1068.230 1433.590 1069.410 1434.770 ;
        RECT 1066.630 1431.990 1067.810 1433.170 ;
        RECT 1068.230 1431.990 1069.410 1433.170 ;
        RECT 1066.630 1253.590 1067.810 1254.770 ;
        RECT 1068.230 1253.590 1069.410 1254.770 ;
        RECT 1066.630 1251.990 1067.810 1253.170 ;
        RECT 1068.230 1251.990 1069.410 1253.170 ;
        RECT 1066.630 1073.590 1067.810 1074.770 ;
        RECT 1068.230 1073.590 1069.410 1074.770 ;
        RECT 1066.630 1071.990 1067.810 1073.170 ;
        RECT 1068.230 1071.990 1069.410 1073.170 ;
        RECT 1066.630 893.590 1067.810 894.770 ;
        RECT 1068.230 893.590 1069.410 894.770 ;
        RECT 1066.630 891.990 1067.810 893.170 ;
        RECT 1068.230 891.990 1069.410 893.170 ;
        RECT 1066.630 713.590 1067.810 714.770 ;
        RECT 1068.230 713.590 1069.410 714.770 ;
        RECT 1066.630 711.990 1067.810 713.170 ;
        RECT 1068.230 711.990 1069.410 713.170 ;
        RECT 1066.630 533.590 1067.810 534.770 ;
        RECT 1068.230 533.590 1069.410 534.770 ;
        RECT 1066.630 531.990 1067.810 533.170 ;
        RECT 1068.230 531.990 1069.410 533.170 ;
        RECT 1066.630 353.590 1067.810 354.770 ;
        RECT 1068.230 353.590 1069.410 354.770 ;
        RECT 1066.630 351.990 1067.810 353.170 ;
        RECT 1068.230 351.990 1069.410 353.170 ;
        RECT 1066.630 173.590 1067.810 174.770 ;
        RECT 1068.230 173.590 1069.410 174.770 ;
        RECT 1066.630 171.990 1067.810 173.170 ;
        RECT 1068.230 171.990 1069.410 173.170 ;
        RECT 1066.630 -36.510 1067.810 -35.330 ;
        RECT 1068.230 -36.510 1069.410 -35.330 ;
        RECT 1066.630 -38.110 1067.810 -36.930 ;
        RECT 1068.230 -38.110 1069.410 -36.930 ;
        RECT 1246.630 3556.610 1247.810 3557.790 ;
        RECT 1248.230 3556.610 1249.410 3557.790 ;
        RECT 1246.630 3555.010 1247.810 3556.190 ;
        RECT 1248.230 3555.010 1249.410 3556.190 ;
        RECT 1246.630 3413.590 1247.810 3414.770 ;
        RECT 1248.230 3413.590 1249.410 3414.770 ;
        RECT 1246.630 3411.990 1247.810 3413.170 ;
        RECT 1248.230 3411.990 1249.410 3413.170 ;
        RECT 1246.630 3233.590 1247.810 3234.770 ;
        RECT 1248.230 3233.590 1249.410 3234.770 ;
        RECT 1246.630 3231.990 1247.810 3233.170 ;
        RECT 1248.230 3231.990 1249.410 3233.170 ;
        RECT 1246.630 3053.590 1247.810 3054.770 ;
        RECT 1248.230 3053.590 1249.410 3054.770 ;
        RECT 1246.630 3051.990 1247.810 3053.170 ;
        RECT 1248.230 3051.990 1249.410 3053.170 ;
        RECT 1246.630 2873.590 1247.810 2874.770 ;
        RECT 1248.230 2873.590 1249.410 2874.770 ;
        RECT 1246.630 2871.990 1247.810 2873.170 ;
        RECT 1248.230 2871.990 1249.410 2873.170 ;
        RECT 1246.630 2693.590 1247.810 2694.770 ;
        RECT 1248.230 2693.590 1249.410 2694.770 ;
        RECT 1246.630 2691.990 1247.810 2693.170 ;
        RECT 1248.230 2691.990 1249.410 2693.170 ;
        RECT 1246.630 2513.590 1247.810 2514.770 ;
        RECT 1248.230 2513.590 1249.410 2514.770 ;
        RECT 1246.630 2511.990 1247.810 2513.170 ;
        RECT 1248.230 2511.990 1249.410 2513.170 ;
        RECT 1246.630 2333.590 1247.810 2334.770 ;
        RECT 1248.230 2333.590 1249.410 2334.770 ;
        RECT 1246.630 2331.990 1247.810 2333.170 ;
        RECT 1248.230 2331.990 1249.410 2333.170 ;
        RECT 1246.630 2153.590 1247.810 2154.770 ;
        RECT 1248.230 2153.590 1249.410 2154.770 ;
        RECT 1246.630 2151.990 1247.810 2153.170 ;
        RECT 1248.230 2151.990 1249.410 2153.170 ;
        RECT 1246.630 1973.590 1247.810 1974.770 ;
        RECT 1248.230 1973.590 1249.410 1974.770 ;
        RECT 1246.630 1971.990 1247.810 1973.170 ;
        RECT 1248.230 1971.990 1249.410 1973.170 ;
        RECT 1246.630 1793.590 1247.810 1794.770 ;
        RECT 1248.230 1793.590 1249.410 1794.770 ;
        RECT 1246.630 1791.990 1247.810 1793.170 ;
        RECT 1248.230 1791.990 1249.410 1793.170 ;
        RECT 1246.630 1613.590 1247.810 1614.770 ;
        RECT 1248.230 1613.590 1249.410 1614.770 ;
        RECT 1246.630 1611.990 1247.810 1613.170 ;
        RECT 1248.230 1611.990 1249.410 1613.170 ;
        RECT 1246.630 1433.590 1247.810 1434.770 ;
        RECT 1248.230 1433.590 1249.410 1434.770 ;
        RECT 1246.630 1431.990 1247.810 1433.170 ;
        RECT 1248.230 1431.990 1249.410 1433.170 ;
        RECT 1246.630 1253.590 1247.810 1254.770 ;
        RECT 1248.230 1253.590 1249.410 1254.770 ;
        RECT 1246.630 1251.990 1247.810 1253.170 ;
        RECT 1248.230 1251.990 1249.410 1253.170 ;
        RECT 1246.630 1073.590 1247.810 1074.770 ;
        RECT 1248.230 1073.590 1249.410 1074.770 ;
        RECT 1246.630 1071.990 1247.810 1073.170 ;
        RECT 1248.230 1071.990 1249.410 1073.170 ;
        RECT 1246.630 893.590 1247.810 894.770 ;
        RECT 1248.230 893.590 1249.410 894.770 ;
        RECT 1246.630 891.990 1247.810 893.170 ;
        RECT 1248.230 891.990 1249.410 893.170 ;
        RECT 1246.630 713.590 1247.810 714.770 ;
        RECT 1248.230 713.590 1249.410 714.770 ;
        RECT 1246.630 711.990 1247.810 713.170 ;
        RECT 1248.230 711.990 1249.410 713.170 ;
        RECT 1246.630 533.590 1247.810 534.770 ;
        RECT 1248.230 533.590 1249.410 534.770 ;
        RECT 1246.630 531.990 1247.810 533.170 ;
        RECT 1248.230 531.990 1249.410 533.170 ;
        RECT 1246.630 353.590 1247.810 354.770 ;
        RECT 1248.230 353.590 1249.410 354.770 ;
        RECT 1246.630 351.990 1247.810 353.170 ;
        RECT 1248.230 351.990 1249.410 353.170 ;
        RECT 1246.630 173.590 1247.810 174.770 ;
        RECT 1248.230 173.590 1249.410 174.770 ;
        RECT 1246.630 171.990 1247.810 173.170 ;
        RECT 1248.230 171.990 1249.410 173.170 ;
        RECT 1246.630 -36.510 1247.810 -35.330 ;
        RECT 1248.230 -36.510 1249.410 -35.330 ;
        RECT 1246.630 -38.110 1247.810 -36.930 ;
        RECT 1248.230 -38.110 1249.410 -36.930 ;
        RECT 1426.630 3556.610 1427.810 3557.790 ;
        RECT 1428.230 3556.610 1429.410 3557.790 ;
        RECT 1426.630 3555.010 1427.810 3556.190 ;
        RECT 1428.230 3555.010 1429.410 3556.190 ;
        RECT 1426.630 3413.590 1427.810 3414.770 ;
        RECT 1428.230 3413.590 1429.410 3414.770 ;
        RECT 1426.630 3411.990 1427.810 3413.170 ;
        RECT 1428.230 3411.990 1429.410 3413.170 ;
        RECT 1426.630 3233.590 1427.810 3234.770 ;
        RECT 1428.230 3233.590 1429.410 3234.770 ;
        RECT 1426.630 3231.990 1427.810 3233.170 ;
        RECT 1428.230 3231.990 1429.410 3233.170 ;
        RECT 1426.630 3053.590 1427.810 3054.770 ;
        RECT 1428.230 3053.590 1429.410 3054.770 ;
        RECT 1426.630 3051.990 1427.810 3053.170 ;
        RECT 1428.230 3051.990 1429.410 3053.170 ;
        RECT 1426.630 2873.590 1427.810 2874.770 ;
        RECT 1428.230 2873.590 1429.410 2874.770 ;
        RECT 1426.630 2871.990 1427.810 2873.170 ;
        RECT 1428.230 2871.990 1429.410 2873.170 ;
        RECT 1426.630 2693.590 1427.810 2694.770 ;
        RECT 1428.230 2693.590 1429.410 2694.770 ;
        RECT 1426.630 2691.990 1427.810 2693.170 ;
        RECT 1428.230 2691.990 1429.410 2693.170 ;
        RECT 1426.630 2513.590 1427.810 2514.770 ;
        RECT 1428.230 2513.590 1429.410 2514.770 ;
        RECT 1426.630 2511.990 1427.810 2513.170 ;
        RECT 1428.230 2511.990 1429.410 2513.170 ;
        RECT 1426.630 2333.590 1427.810 2334.770 ;
        RECT 1428.230 2333.590 1429.410 2334.770 ;
        RECT 1426.630 2331.990 1427.810 2333.170 ;
        RECT 1428.230 2331.990 1429.410 2333.170 ;
        RECT 1426.630 2153.590 1427.810 2154.770 ;
        RECT 1428.230 2153.590 1429.410 2154.770 ;
        RECT 1426.630 2151.990 1427.810 2153.170 ;
        RECT 1428.230 2151.990 1429.410 2153.170 ;
        RECT 1426.630 1973.590 1427.810 1974.770 ;
        RECT 1428.230 1973.590 1429.410 1974.770 ;
        RECT 1426.630 1971.990 1427.810 1973.170 ;
        RECT 1428.230 1971.990 1429.410 1973.170 ;
        RECT 1426.630 1793.590 1427.810 1794.770 ;
        RECT 1428.230 1793.590 1429.410 1794.770 ;
        RECT 1426.630 1791.990 1427.810 1793.170 ;
        RECT 1428.230 1791.990 1429.410 1793.170 ;
        RECT 1426.630 1613.590 1427.810 1614.770 ;
        RECT 1428.230 1613.590 1429.410 1614.770 ;
        RECT 1426.630 1611.990 1427.810 1613.170 ;
        RECT 1428.230 1611.990 1429.410 1613.170 ;
        RECT 1426.630 1433.590 1427.810 1434.770 ;
        RECT 1428.230 1433.590 1429.410 1434.770 ;
        RECT 1426.630 1431.990 1427.810 1433.170 ;
        RECT 1428.230 1431.990 1429.410 1433.170 ;
        RECT 1426.630 1253.590 1427.810 1254.770 ;
        RECT 1428.230 1253.590 1429.410 1254.770 ;
        RECT 1426.630 1251.990 1427.810 1253.170 ;
        RECT 1428.230 1251.990 1429.410 1253.170 ;
        RECT 1426.630 1073.590 1427.810 1074.770 ;
        RECT 1428.230 1073.590 1429.410 1074.770 ;
        RECT 1426.630 1071.990 1427.810 1073.170 ;
        RECT 1428.230 1071.990 1429.410 1073.170 ;
        RECT 1426.630 893.590 1427.810 894.770 ;
        RECT 1428.230 893.590 1429.410 894.770 ;
        RECT 1426.630 891.990 1427.810 893.170 ;
        RECT 1428.230 891.990 1429.410 893.170 ;
        RECT 1426.630 713.590 1427.810 714.770 ;
        RECT 1428.230 713.590 1429.410 714.770 ;
        RECT 1426.630 711.990 1427.810 713.170 ;
        RECT 1428.230 711.990 1429.410 713.170 ;
        RECT 1426.630 533.590 1427.810 534.770 ;
        RECT 1428.230 533.590 1429.410 534.770 ;
        RECT 1426.630 531.990 1427.810 533.170 ;
        RECT 1428.230 531.990 1429.410 533.170 ;
        RECT 1426.630 353.590 1427.810 354.770 ;
        RECT 1428.230 353.590 1429.410 354.770 ;
        RECT 1426.630 351.990 1427.810 353.170 ;
        RECT 1428.230 351.990 1429.410 353.170 ;
        RECT 1426.630 173.590 1427.810 174.770 ;
        RECT 1428.230 173.590 1429.410 174.770 ;
        RECT 1426.630 171.990 1427.810 173.170 ;
        RECT 1428.230 171.990 1429.410 173.170 ;
        RECT 1426.630 -36.510 1427.810 -35.330 ;
        RECT 1428.230 -36.510 1429.410 -35.330 ;
        RECT 1426.630 -38.110 1427.810 -36.930 ;
        RECT 1428.230 -38.110 1429.410 -36.930 ;
        RECT 1606.630 3556.610 1607.810 3557.790 ;
        RECT 1608.230 3556.610 1609.410 3557.790 ;
        RECT 1606.630 3555.010 1607.810 3556.190 ;
        RECT 1608.230 3555.010 1609.410 3556.190 ;
        RECT 1606.630 3413.590 1607.810 3414.770 ;
        RECT 1608.230 3413.590 1609.410 3414.770 ;
        RECT 1606.630 3411.990 1607.810 3413.170 ;
        RECT 1608.230 3411.990 1609.410 3413.170 ;
        RECT 1606.630 3233.590 1607.810 3234.770 ;
        RECT 1608.230 3233.590 1609.410 3234.770 ;
        RECT 1606.630 3231.990 1607.810 3233.170 ;
        RECT 1608.230 3231.990 1609.410 3233.170 ;
        RECT 1606.630 3053.590 1607.810 3054.770 ;
        RECT 1608.230 3053.590 1609.410 3054.770 ;
        RECT 1606.630 3051.990 1607.810 3053.170 ;
        RECT 1608.230 3051.990 1609.410 3053.170 ;
        RECT 1606.630 2873.590 1607.810 2874.770 ;
        RECT 1608.230 2873.590 1609.410 2874.770 ;
        RECT 1606.630 2871.990 1607.810 2873.170 ;
        RECT 1608.230 2871.990 1609.410 2873.170 ;
        RECT 1606.630 2693.590 1607.810 2694.770 ;
        RECT 1608.230 2693.590 1609.410 2694.770 ;
        RECT 1606.630 2691.990 1607.810 2693.170 ;
        RECT 1608.230 2691.990 1609.410 2693.170 ;
        RECT 1606.630 2513.590 1607.810 2514.770 ;
        RECT 1608.230 2513.590 1609.410 2514.770 ;
        RECT 1606.630 2511.990 1607.810 2513.170 ;
        RECT 1608.230 2511.990 1609.410 2513.170 ;
        RECT 1606.630 2333.590 1607.810 2334.770 ;
        RECT 1608.230 2333.590 1609.410 2334.770 ;
        RECT 1606.630 2331.990 1607.810 2333.170 ;
        RECT 1608.230 2331.990 1609.410 2333.170 ;
        RECT 1606.630 2153.590 1607.810 2154.770 ;
        RECT 1608.230 2153.590 1609.410 2154.770 ;
        RECT 1606.630 2151.990 1607.810 2153.170 ;
        RECT 1608.230 2151.990 1609.410 2153.170 ;
        RECT 1606.630 1973.590 1607.810 1974.770 ;
        RECT 1608.230 1973.590 1609.410 1974.770 ;
        RECT 1606.630 1971.990 1607.810 1973.170 ;
        RECT 1608.230 1971.990 1609.410 1973.170 ;
        RECT 1606.630 1793.590 1607.810 1794.770 ;
        RECT 1608.230 1793.590 1609.410 1794.770 ;
        RECT 1606.630 1791.990 1607.810 1793.170 ;
        RECT 1608.230 1791.990 1609.410 1793.170 ;
        RECT 1606.630 1613.590 1607.810 1614.770 ;
        RECT 1608.230 1613.590 1609.410 1614.770 ;
        RECT 1606.630 1611.990 1607.810 1613.170 ;
        RECT 1608.230 1611.990 1609.410 1613.170 ;
        RECT 1606.630 1433.590 1607.810 1434.770 ;
        RECT 1608.230 1433.590 1609.410 1434.770 ;
        RECT 1606.630 1431.990 1607.810 1433.170 ;
        RECT 1608.230 1431.990 1609.410 1433.170 ;
        RECT 1606.630 1253.590 1607.810 1254.770 ;
        RECT 1608.230 1253.590 1609.410 1254.770 ;
        RECT 1606.630 1251.990 1607.810 1253.170 ;
        RECT 1608.230 1251.990 1609.410 1253.170 ;
        RECT 1606.630 1073.590 1607.810 1074.770 ;
        RECT 1608.230 1073.590 1609.410 1074.770 ;
        RECT 1606.630 1071.990 1607.810 1073.170 ;
        RECT 1608.230 1071.990 1609.410 1073.170 ;
        RECT 1606.630 893.590 1607.810 894.770 ;
        RECT 1608.230 893.590 1609.410 894.770 ;
        RECT 1606.630 891.990 1607.810 893.170 ;
        RECT 1608.230 891.990 1609.410 893.170 ;
        RECT 1606.630 713.590 1607.810 714.770 ;
        RECT 1608.230 713.590 1609.410 714.770 ;
        RECT 1606.630 711.990 1607.810 713.170 ;
        RECT 1608.230 711.990 1609.410 713.170 ;
        RECT 1606.630 533.590 1607.810 534.770 ;
        RECT 1608.230 533.590 1609.410 534.770 ;
        RECT 1606.630 531.990 1607.810 533.170 ;
        RECT 1608.230 531.990 1609.410 533.170 ;
        RECT 1606.630 353.590 1607.810 354.770 ;
        RECT 1608.230 353.590 1609.410 354.770 ;
        RECT 1606.630 351.990 1607.810 353.170 ;
        RECT 1608.230 351.990 1609.410 353.170 ;
        RECT 1606.630 173.590 1607.810 174.770 ;
        RECT 1608.230 173.590 1609.410 174.770 ;
        RECT 1606.630 171.990 1607.810 173.170 ;
        RECT 1608.230 171.990 1609.410 173.170 ;
        RECT 1606.630 -36.510 1607.810 -35.330 ;
        RECT 1608.230 -36.510 1609.410 -35.330 ;
        RECT 1606.630 -38.110 1607.810 -36.930 ;
        RECT 1608.230 -38.110 1609.410 -36.930 ;
        RECT 1786.630 3556.610 1787.810 3557.790 ;
        RECT 1788.230 3556.610 1789.410 3557.790 ;
        RECT 1786.630 3555.010 1787.810 3556.190 ;
        RECT 1788.230 3555.010 1789.410 3556.190 ;
        RECT 1786.630 3413.590 1787.810 3414.770 ;
        RECT 1788.230 3413.590 1789.410 3414.770 ;
        RECT 1786.630 3411.990 1787.810 3413.170 ;
        RECT 1788.230 3411.990 1789.410 3413.170 ;
        RECT 1786.630 3233.590 1787.810 3234.770 ;
        RECT 1788.230 3233.590 1789.410 3234.770 ;
        RECT 1786.630 3231.990 1787.810 3233.170 ;
        RECT 1788.230 3231.990 1789.410 3233.170 ;
        RECT 1786.630 3053.590 1787.810 3054.770 ;
        RECT 1788.230 3053.590 1789.410 3054.770 ;
        RECT 1786.630 3051.990 1787.810 3053.170 ;
        RECT 1788.230 3051.990 1789.410 3053.170 ;
        RECT 1786.630 2873.590 1787.810 2874.770 ;
        RECT 1788.230 2873.590 1789.410 2874.770 ;
        RECT 1786.630 2871.990 1787.810 2873.170 ;
        RECT 1788.230 2871.990 1789.410 2873.170 ;
        RECT 1786.630 2693.590 1787.810 2694.770 ;
        RECT 1788.230 2693.590 1789.410 2694.770 ;
        RECT 1786.630 2691.990 1787.810 2693.170 ;
        RECT 1788.230 2691.990 1789.410 2693.170 ;
        RECT 1786.630 2513.590 1787.810 2514.770 ;
        RECT 1788.230 2513.590 1789.410 2514.770 ;
        RECT 1786.630 2511.990 1787.810 2513.170 ;
        RECT 1788.230 2511.990 1789.410 2513.170 ;
        RECT 1786.630 2333.590 1787.810 2334.770 ;
        RECT 1788.230 2333.590 1789.410 2334.770 ;
        RECT 1786.630 2331.990 1787.810 2333.170 ;
        RECT 1788.230 2331.990 1789.410 2333.170 ;
        RECT 1786.630 2153.590 1787.810 2154.770 ;
        RECT 1788.230 2153.590 1789.410 2154.770 ;
        RECT 1786.630 2151.990 1787.810 2153.170 ;
        RECT 1788.230 2151.990 1789.410 2153.170 ;
        RECT 1786.630 1973.590 1787.810 1974.770 ;
        RECT 1788.230 1973.590 1789.410 1974.770 ;
        RECT 1786.630 1971.990 1787.810 1973.170 ;
        RECT 1788.230 1971.990 1789.410 1973.170 ;
        RECT 1786.630 1793.590 1787.810 1794.770 ;
        RECT 1788.230 1793.590 1789.410 1794.770 ;
        RECT 1786.630 1791.990 1787.810 1793.170 ;
        RECT 1788.230 1791.990 1789.410 1793.170 ;
        RECT 1786.630 1613.590 1787.810 1614.770 ;
        RECT 1788.230 1613.590 1789.410 1614.770 ;
        RECT 1786.630 1611.990 1787.810 1613.170 ;
        RECT 1788.230 1611.990 1789.410 1613.170 ;
        RECT 1786.630 1433.590 1787.810 1434.770 ;
        RECT 1788.230 1433.590 1789.410 1434.770 ;
        RECT 1786.630 1431.990 1787.810 1433.170 ;
        RECT 1788.230 1431.990 1789.410 1433.170 ;
        RECT 1786.630 1253.590 1787.810 1254.770 ;
        RECT 1788.230 1253.590 1789.410 1254.770 ;
        RECT 1786.630 1251.990 1787.810 1253.170 ;
        RECT 1788.230 1251.990 1789.410 1253.170 ;
        RECT 1786.630 1073.590 1787.810 1074.770 ;
        RECT 1788.230 1073.590 1789.410 1074.770 ;
        RECT 1786.630 1071.990 1787.810 1073.170 ;
        RECT 1788.230 1071.990 1789.410 1073.170 ;
        RECT 1786.630 893.590 1787.810 894.770 ;
        RECT 1788.230 893.590 1789.410 894.770 ;
        RECT 1786.630 891.990 1787.810 893.170 ;
        RECT 1788.230 891.990 1789.410 893.170 ;
        RECT 1786.630 713.590 1787.810 714.770 ;
        RECT 1788.230 713.590 1789.410 714.770 ;
        RECT 1786.630 711.990 1787.810 713.170 ;
        RECT 1788.230 711.990 1789.410 713.170 ;
        RECT 1786.630 533.590 1787.810 534.770 ;
        RECT 1788.230 533.590 1789.410 534.770 ;
        RECT 1786.630 531.990 1787.810 533.170 ;
        RECT 1788.230 531.990 1789.410 533.170 ;
        RECT 1786.630 353.590 1787.810 354.770 ;
        RECT 1788.230 353.590 1789.410 354.770 ;
        RECT 1786.630 351.990 1787.810 353.170 ;
        RECT 1788.230 351.990 1789.410 353.170 ;
        RECT 1786.630 173.590 1787.810 174.770 ;
        RECT 1788.230 173.590 1789.410 174.770 ;
        RECT 1786.630 171.990 1787.810 173.170 ;
        RECT 1788.230 171.990 1789.410 173.170 ;
        RECT 1786.630 -36.510 1787.810 -35.330 ;
        RECT 1788.230 -36.510 1789.410 -35.330 ;
        RECT 1786.630 -38.110 1787.810 -36.930 ;
        RECT 1788.230 -38.110 1789.410 -36.930 ;
        RECT 1966.630 3556.610 1967.810 3557.790 ;
        RECT 1968.230 3556.610 1969.410 3557.790 ;
        RECT 1966.630 3555.010 1967.810 3556.190 ;
        RECT 1968.230 3555.010 1969.410 3556.190 ;
        RECT 1966.630 3413.590 1967.810 3414.770 ;
        RECT 1968.230 3413.590 1969.410 3414.770 ;
        RECT 1966.630 3411.990 1967.810 3413.170 ;
        RECT 1968.230 3411.990 1969.410 3413.170 ;
        RECT 1966.630 3233.590 1967.810 3234.770 ;
        RECT 1968.230 3233.590 1969.410 3234.770 ;
        RECT 1966.630 3231.990 1967.810 3233.170 ;
        RECT 1968.230 3231.990 1969.410 3233.170 ;
        RECT 1966.630 3053.590 1967.810 3054.770 ;
        RECT 1968.230 3053.590 1969.410 3054.770 ;
        RECT 1966.630 3051.990 1967.810 3053.170 ;
        RECT 1968.230 3051.990 1969.410 3053.170 ;
        RECT 1966.630 2873.590 1967.810 2874.770 ;
        RECT 1968.230 2873.590 1969.410 2874.770 ;
        RECT 1966.630 2871.990 1967.810 2873.170 ;
        RECT 1968.230 2871.990 1969.410 2873.170 ;
        RECT 1966.630 2693.590 1967.810 2694.770 ;
        RECT 1968.230 2693.590 1969.410 2694.770 ;
        RECT 1966.630 2691.990 1967.810 2693.170 ;
        RECT 1968.230 2691.990 1969.410 2693.170 ;
        RECT 1966.630 2513.590 1967.810 2514.770 ;
        RECT 1968.230 2513.590 1969.410 2514.770 ;
        RECT 1966.630 2511.990 1967.810 2513.170 ;
        RECT 1968.230 2511.990 1969.410 2513.170 ;
        RECT 1966.630 2333.590 1967.810 2334.770 ;
        RECT 1968.230 2333.590 1969.410 2334.770 ;
        RECT 1966.630 2331.990 1967.810 2333.170 ;
        RECT 1968.230 2331.990 1969.410 2333.170 ;
        RECT 1966.630 2153.590 1967.810 2154.770 ;
        RECT 1968.230 2153.590 1969.410 2154.770 ;
        RECT 1966.630 2151.990 1967.810 2153.170 ;
        RECT 1968.230 2151.990 1969.410 2153.170 ;
        RECT 1966.630 1973.590 1967.810 1974.770 ;
        RECT 1968.230 1973.590 1969.410 1974.770 ;
        RECT 1966.630 1971.990 1967.810 1973.170 ;
        RECT 1968.230 1971.990 1969.410 1973.170 ;
        RECT 1966.630 1793.590 1967.810 1794.770 ;
        RECT 1968.230 1793.590 1969.410 1794.770 ;
        RECT 1966.630 1791.990 1967.810 1793.170 ;
        RECT 1968.230 1791.990 1969.410 1793.170 ;
        RECT 1966.630 1613.590 1967.810 1614.770 ;
        RECT 1968.230 1613.590 1969.410 1614.770 ;
        RECT 1966.630 1611.990 1967.810 1613.170 ;
        RECT 1968.230 1611.990 1969.410 1613.170 ;
        RECT 1966.630 1433.590 1967.810 1434.770 ;
        RECT 1968.230 1433.590 1969.410 1434.770 ;
        RECT 1966.630 1431.990 1967.810 1433.170 ;
        RECT 1968.230 1431.990 1969.410 1433.170 ;
        RECT 1966.630 1253.590 1967.810 1254.770 ;
        RECT 1968.230 1253.590 1969.410 1254.770 ;
        RECT 1966.630 1251.990 1967.810 1253.170 ;
        RECT 1968.230 1251.990 1969.410 1253.170 ;
        RECT 1966.630 1073.590 1967.810 1074.770 ;
        RECT 1968.230 1073.590 1969.410 1074.770 ;
        RECT 1966.630 1071.990 1967.810 1073.170 ;
        RECT 1968.230 1071.990 1969.410 1073.170 ;
        RECT 1966.630 893.590 1967.810 894.770 ;
        RECT 1968.230 893.590 1969.410 894.770 ;
        RECT 1966.630 891.990 1967.810 893.170 ;
        RECT 1968.230 891.990 1969.410 893.170 ;
        RECT 1966.630 713.590 1967.810 714.770 ;
        RECT 1968.230 713.590 1969.410 714.770 ;
        RECT 1966.630 711.990 1967.810 713.170 ;
        RECT 1968.230 711.990 1969.410 713.170 ;
        RECT 1966.630 533.590 1967.810 534.770 ;
        RECT 1968.230 533.590 1969.410 534.770 ;
        RECT 1966.630 531.990 1967.810 533.170 ;
        RECT 1968.230 531.990 1969.410 533.170 ;
        RECT 1966.630 353.590 1967.810 354.770 ;
        RECT 1968.230 353.590 1969.410 354.770 ;
        RECT 1966.630 351.990 1967.810 353.170 ;
        RECT 1968.230 351.990 1969.410 353.170 ;
        RECT 1966.630 173.590 1967.810 174.770 ;
        RECT 1968.230 173.590 1969.410 174.770 ;
        RECT 1966.630 171.990 1967.810 173.170 ;
        RECT 1968.230 171.990 1969.410 173.170 ;
        RECT 1966.630 -36.510 1967.810 -35.330 ;
        RECT 1968.230 -36.510 1969.410 -35.330 ;
        RECT 1966.630 -38.110 1967.810 -36.930 ;
        RECT 1968.230 -38.110 1969.410 -36.930 ;
        RECT 2146.630 3556.610 2147.810 3557.790 ;
        RECT 2148.230 3556.610 2149.410 3557.790 ;
        RECT 2146.630 3555.010 2147.810 3556.190 ;
        RECT 2148.230 3555.010 2149.410 3556.190 ;
        RECT 2146.630 3413.590 2147.810 3414.770 ;
        RECT 2148.230 3413.590 2149.410 3414.770 ;
        RECT 2146.630 3411.990 2147.810 3413.170 ;
        RECT 2148.230 3411.990 2149.410 3413.170 ;
        RECT 2146.630 3233.590 2147.810 3234.770 ;
        RECT 2148.230 3233.590 2149.410 3234.770 ;
        RECT 2146.630 3231.990 2147.810 3233.170 ;
        RECT 2148.230 3231.990 2149.410 3233.170 ;
        RECT 2146.630 3053.590 2147.810 3054.770 ;
        RECT 2148.230 3053.590 2149.410 3054.770 ;
        RECT 2146.630 3051.990 2147.810 3053.170 ;
        RECT 2148.230 3051.990 2149.410 3053.170 ;
        RECT 2146.630 2873.590 2147.810 2874.770 ;
        RECT 2148.230 2873.590 2149.410 2874.770 ;
        RECT 2146.630 2871.990 2147.810 2873.170 ;
        RECT 2148.230 2871.990 2149.410 2873.170 ;
        RECT 2146.630 2693.590 2147.810 2694.770 ;
        RECT 2148.230 2693.590 2149.410 2694.770 ;
        RECT 2146.630 2691.990 2147.810 2693.170 ;
        RECT 2148.230 2691.990 2149.410 2693.170 ;
        RECT 2146.630 2513.590 2147.810 2514.770 ;
        RECT 2148.230 2513.590 2149.410 2514.770 ;
        RECT 2146.630 2511.990 2147.810 2513.170 ;
        RECT 2148.230 2511.990 2149.410 2513.170 ;
        RECT 2146.630 2333.590 2147.810 2334.770 ;
        RECT 2148.230 2333.590 2149.410 2334.770 ;
        RECT 2146.630 2331.990 2147.810 2333.170 ;
        RECT 2148.230 2331.990 2149.410 2333.170 ;
        RECT 2146.630 2153.590 2147.810 2154.770 ;
        RECT 2148.230 2153.590 2149.410 2154.770 ;
        RECT 2146.630 2151.990 2147.810 2153.170 ;
        RECT 2148.230 2151.990 2149.410 2153.170 ;
        RECT 2146.630 1973.590 2147.810 1974.770 ;
        RECT 2148.230 1973.590 2149.410 1974.770 ;
        RECT 2146.630 1971.990 2147.810 1973.170 ;
        RECT 2148.230 1971.990 2149.410 1973.170 ;
        RECT 2146.630 1793.590 2147.810 1794.770 ;
        RECT 2148.230 1793.590 2149.410 1794.770 ;
        RECT 2146.630 1791.990 2147.810 1793.170 ;
        RECT 2148.230 1791.990 2149.410 1793.170 ;
        RECT 2146.630 1613.590 2147.810 1614.770 ;
        RECT 2148.230 1613.590 2149.410 1614.770 ;
        RECT 2146.630 1611.990 2147.810 1613.170 ;
        RECT 2148.230 1611.990 2149.410 1613.170 ;
        RECT 2146.630 1433.590 2147.810 1434.770 ;
        RECT 2148.230 1433.590 2149.410 1434.770 ;
        RECT 2146.630 1431.990 2147.810 1433.170 ;
        RECT 2148.230 1431.990 2149.410 1433.170 ;
        RECT 2146.630 1253.590 2147.810 1254.770 ;
        RECT 2148.230 1253.590 2149.410 1254.770 ;
        RECT 2146.630 1251.990 2147.810 1253.170 ;
        RECT 2148.230 1251.990 2149.410 1253.170 ;
        RECT 2146.630 1073.590 2147.810 1074.770 ;
        RECT 2148.230 1073.590 2149.410 1074.770 ;
        RECT 2146.630 1071.990 2147.810 1073.170 ;
        RECT 2148.230 1071.990 2149.410 1073.170 ;
        RECT 2146.630 893.590 2147.810 894.770 ;
        RECT 2148.230 893.590 2149.410 894.770 ;
        RECT 2146.630 891.990 2147.810 893.170 ;
        RECT 2148.230 891.990 2149.410 893.170 ;
        RECT 2146.630 713.590 2147.810 714.770 ;
        RECT 2148.230 713.590 2149.410 714.770 ;
        RECT 2146.630 711.990 2147.810 713.170 ;
        RECT 2148.230 711.990 2149.410 713.170 ;
        RECT 2146.630 533.590 2147.810 534.770 ;
        RECT 2148.230 533.590 2149.410 534.770 ;
        RECT 2146.630 531.990 2147.810 533.170 ;
        RECT 2148.230 531.990 2149.410 533.170 ;
        RECT 2146.630 353.590 2147.810 354.770 ;
        RECT 2148.230 353.590 2149.410 354.770 ;
        RECT 2146.630 351.990 2147.810 353.170 ;
        RECT 2148.230 351.990 2149.410 353.170 ;
        RECT 2146.630 173.590 2147.810 174.770 ;
        RECT 2148.230 173.590 2149.410 174.770 ;
        RECT 2146.630 171.990 2147.810 173.170 ;
        RECT 2148.230 171.990 2149.410 173.170 ;
        RECT 2146.630 -36.510 2147.810 -35.330 ;
        RECT 2148.230 -36.510 2149.410 -35.330 ;
        RECT 2146.630 -38.110 2147.810 -36.930 ;
        RECT 2148.230 -38.110 2149.410 -36.930 ;
        RECT 2326.630 3556.610 2327.810 3557.790 ;
        RECT 2328.230 3556.610 2329.410 3557.790 ;
        RECT 2326.630 3555.010 2327.810 3556.190 ;
        RECT 2328.230 3555.010 2329.410 3556.190 ;
        RECT 2326.630 3413.590 2327.810 3414.770 ;
        RECT 2328.230 3413.590 2329.410 3414.770 ;
        RECT 2326.630 3411.990 2327.810 3413.170 ;
        RECT 2328.230 3411.990 2329.410 3413.170 ;
        RECT 2326.630 3233.590 2327.810 3234.770 ;
        RECT 2328.230 3233.590 2329.410 3234.770 ;
        RECT 2326.630 3231.990 2327.810 3233.170 ;
        RECT 2328.230 3231.990 2329.410 3233.170 ;
        RECT 2326.630 3053.590 2327.810 3054.770 ;
        RECT 2328.230 3053.590 2329.410 3054.770 ;
        RECT 2326.630 3051.990 2327.810 3053.170 ;
        RECT 2328.230 3051.990 2329.410 3053.170 ;
        RECT 2326.630 2873.590 2327.810 2874.770 ;
        RECT 2328.230 2873.590 2329.410 2874.770 ;
        RECT 2326.630 2871.990 2327.810 2873.170 ;
        RECT 2328.230 2871.990 2329.410 2873.170 ;
        RECT 2326.630 2693.590 2327.810 2694.770 ;
        RECT 2328.230 2693.590 2329.410 2694.770 ;
        RECT 2326.630 2691.990 2327.810 2693.170 ;
        RECT 2328.230 2691.990 2329.410 2693.170 ;
        RECT 2326.630 2513.590 2327.810 2514.770 ;
        RECT 2328.230 2513.590 2329.410 2514.770 ;
        RECT 2326.630 2511.990 2327.810 2513.170 ;
        RECT 2328.230 2511.990 2329.410 2513.170 ;
        RECT 2326.630 2333.590 2327.810 2334.770 ;
        RECT 2328.230 2333.590 2329.410 2334.770 ;
        RECT 2326.630 2331.990 2327.810 2333.170 ;
        RECT 2328.230 2331.990 2329.410 2333.170 ;
        RECT 2326.630 2153.590 2327.810 2154.770 ;
        RECT 2328.230 2153.590 2329.410 2154.770 ;
        RECT 2326.630 2151.990 2327.810 2153.170 ;
        RECT 2328.230 2151.990 2329.410 2153.170 ;
        RECT 2326.630 1973.590 2327.810 1974.770 ;
        RECT 2328.230 1973.590 2329.410 1974.770 ;
        RECT 2326.630 1971.990 2327.810 1973.170 ;
        RECT 2328.230 1971.990 2329.410 1973.170 ;
        RECT 2326.630 1793.590 2327.810 1794.770 ;
        RECT 2328.230 1793.590 2329.410 1794.770 ;
        RECT 2326.630 1791.990 2327.810 1793.170 ;
        RECT 2328.230 1791.990 2329.410 1793.170 ;
        RECT 2326.630 1613.590 2327.810 1614.770 ;
        RECT 2328.230 1613.590 2329.410 1614.770 ;
        RECT 2326.630 1611.990 2327.810 1613.170 ;
        RECT 2328.230 1611.990 2329.410 1613.170 ;
        RECT 2326.630 1433.590 2327.810 1434.770 ;
        RECT 2328.230 1433.590 2329.410 1434.770 ;
        RECT 2326.630 1431.990 2327.810 1433.170 ;
        RECT 2328.230 1431.990 2329.410 1433.170 ;
        RECT 2326.630 1253.590 2327.810 1254.770 ;
        RECT 2328.230 1253.590 2329.410 1254.770 ;
        RECT 2326.630 1251.990 2327.810 1253.170 ;
        RECT 2328.230 1251.990 2329.410 1253.170 ;
        RECT 2326.630 1073.590 2327.810 1074.770 ;
        RECT 2328.230 1073.590 2329.410 1074.770 ;
        RECT 2326.630 1071.990 2327.810 1073.170 ;
        RECT 2328.230 1071.990 2329.410 1073.170 ;
        RECT 2326.630 893.590 2327.810 894.770 ;
        RECT 2328.230 893.590 2329.410 894.770 ;
        RECT 2326.630 891.990 2327.810 893.170 ;
        RECT 2328.230 891.990 2329.410 893.170 ;
        RECT 2326.630 713.590 2327.810 714.770 ;
        RECT 2328.230 713.590 2329.410 714.770 ;
        RECT 2326.630 711.990 2327.810 713.170 ;
        RECT 2328.230 711.990 2329.410 713.170 ;
        RECT 2326.630 533.590 2327.810 534.770 ;
        RECT 2328.230 533.590 2329.410 534.770 ;
        RECT 2326.630 531.990 2327.810 533.170 ;
        RECT 2328.230 531.990 2329.410 533.170 ;
        RECT 2326.630 353.590 2327.810 354.770 ;
        RECT 2328.230 353.590 2329.410 354.770 ;
        RECT 2326.630 351.990 2327.810 353.170 ;
        RECT 2328.230 351.990 2329.410 353.170 ;
        RECT 2326.630 173.590 2327.810 174.770 ;
        RECT 2328.230 173.590 2329.410 174.770 ;
        RECT 2326.630 171.990 2327.810 173.170 ;
        RECT 2328.230 171.990 2329.410 173.170 ;
        RECT 2326.630 -36.510 2327.810 -35.330 ;
        RECT 2328.230 -36.510 2329.410 -35.330 ;
        RECT 2326.630 -38.110 2327.810 -36.930 ;
        RECT 2328.230 -38.110 2329.410 -36.930 ;
        RECT 2506.630 3556.610 2507.810 3557.790 ;
        RECT 2508.230 3556.610 2509.410 3557.790 ;
        RECT 2506.630 3555.010 2507.810 3556.190 ;
        RECT 2508.230 3555.010 2509.410 3556.190 ;
        RECT 2506.630 3413.590 2507.810 3414.770 ;
        RECT 2508.230 3413.590 2509.410 3414.770 ;
        RECT 2506.630 3411.990 2507.810 3413.170 ;
        RECT 2508.230 3411.990 2509.410 3413.170 ;
        RECT 2506.630 3233.590 2507.810 3234.770 ;
        RECT 2508.230 3233.590 2509.410 3234.770 ;
        RECT 2506.630 3231.990 2507.810 3233.170 ;
        RECT 2508.230 3231.990 2509.410 3233.170 ;
        RECT 2506.630 3053.590 2507.810 3054.770 ;
        RECT 2508.230 3053.590 2509.410 3054.770 ;
        RECT 2506.630 3051.990 2507.810 3053.170 ;
        RECT 2508.230 3051.990 2509.410 3053.170 ;
        RECT 2506.630 2873.590 2507.810 2874.770 ;
        RECT 2508.230 2873.590 2509.410 2874.770 ;
        RECT 2506.630 2871.990 2507.810 2873.170 ;
        RECT 2508.230 2871.990 2509.410 2873.170 ;
        RECT 2506.630 2693.590 2507.810 2694.770 ;
        RECT 2508.230 2693.590 2509.410 2694.770 ;
        RECT 2506.630 2691.990 2507.810 2693.170 ;
        RECT 2508.230 2691.990 2509.410 2693.170 ;
        RECT 2506.630 2513.590 2507.810 2514.770 ;
        RECT 2508.230 2513.590 2509.410 2514.770 ;
        RECT 2506.630 2511.990 2507.810 2513.170 ;
        RECT 2508.230 2511.990 2509.410 2513.170 ;
        RECT 2506.630 2333.590 2507.810 2334.770 ;
        RECT 2508.230 2333.590 2509.410 2334.770 ;
        RECT 2506.630 2331.990 2507.810 2333.170 ;
        RECT 2508.230 2331.990 2509.410 2333.170 ;
        RECT 2506.630 2153.590 2507.810 2154.770 ;
        RECT 2508.230 2153.590 2509.410 2154.770 ;
        RECT 2506.630 2151.990 2507.810 2153.170 ;
        RECT 2508.230 2151.990 2509.410 2153.170 ;
        RECT 2506.630 1973.590 2507.810 1974.770 ;
        RECT 2508.230 1973.590 2509.410 1974.770 ;
        RECT 2506.630 1971.990 2507.810 1973.170 ;
        RECT 2508.230 1971.990 2509.410 1973.170 ;
        RECT 2506.630 1793.590 2507.810 1794.770 ;
        RECT 2508.230 1793.590 2509.410 1794.770 ;
        RECT 2506.630 1791.990 2507.810 1793.170 ;
        RECT 2508.230 1791.990 2509.410 1793.170 ;
        RECT 2506.630 1613.590 2507.810 1614.770 ;
        RECT 2508.230 1613.590 2509.410 1614.770 ;
        RECT 2506.630 1611.990 2507.810 1613.170 ;
        RECT 2508.230 1611.990 2509.410 1613.170 ;
        RECT 2506.630 1433.590 2507.810 1434.770 ;
        RECT 2508.230 1433.590 2509.410 1434.770 ;
        RECT 2506.630 1431.990 2507.810 1433.170 ;
        RECT 2508.230 1431.990 2509.410 1433.170 ;
        RECT 2506.630 1253.590 2507.810 1254.770 ;
        RECT 2508.230 1253.590 2509.410 1254.770 ;
        RECT 2506.630 1251.990 2507.810 1253.170 ;
        RECT 2508.230 1251.990 2509.410 1253.170 ;
        RECT 2506.630 1073.590 2507.810 1074.770 ;
        RECT 2508.230 1073.590 2509.410 1074.770 ;
        RECT 2506.630 1071.990 2507.810 1073.170 ;
        RECT 2508.230 1071.990 2509.410 1073.170 ;
        RECT 2506.630 893.590 2507.810 894.770 ;
        RECT 2508.230 893.590 2509.410 894.770 ;
        RECT 2506.630 891.990 2507.810 893.170 ;
        RECT 2508.230 891.990 2509.410 893.170 ;
        RECT 2506.630 713.590 2507.810 714.770 ;
        RECT 2508.230 713.590 2509.410 714.770 ;
        RECT 2506.630 711.990 2507.810 713.170 ;
        RECT 2508.230 711.990 2509.410 713.170 ;
        RECT 2506.630 533.590 2507.810 534.770 ;
        RECT 2508.230 533.590 2509.410 534.770 ;
        RECT 2506.630 531.990 2507.810 533.170 ;
        RECT 2508.230 531.990 2509.410 533.170 ;
        RECT 2506.630 353.590 2507.810 354.770 ;
        RECT 2508.230 353.590 2509.410 354.770 ;
        RECT 2506.630 351.990 2507.810 353.170 ;
        RECT 2508.230 351.990 2509.410 353.170 ;
        RECT 2506.630 173.590 2507.810 174.770 ;
        RECT 2508.230 173.590 2509.410 174.770 ;
        RECT 2506.630 171.990 2507.810 173.170 ;
        RECT 2508.230 171.990 2509.410 173.170 ;
        RECT 2506.630 -36.510 2507.810 -35.330 ;
        RECT 2508.230 -36.510 2509.410 -35.330 ;
        RECT 2506.630 -38.110 2507.810 -36.930 ;
        RECT 2508.230 -38.110 2509.410 -36.930 ;
        RECT 2686.630 3556.610 2687.810 3557.790 ;
        RECT 2688.230 3556.610 2689.410 3557.790 ;
        RECT 2686.630 3555.010 2687.810 3556.190 ;
        RECT 2688.230 3555.010 2689.410 3556.190 ;
        RECT 2686.630 3413.590 2687.810 3414.770 ;
        RECT 2688.230 3413.590 2689.410 3414.770 ;
        RECT 2686.630 3411.990 2687.810 3413.170 ;
        RECT 2688.230 3411.990 2689.410 3413.170 ;
        RECT 2686.630 3233.590 2687.810 3234.770 ;
        RECT 2688.230 3233.590 2689.410 3234.770 ;
        RECT 2686.630 3231.990 2687.810 3233.170 ;
        RECT 2688.230 3231.990 2689.410 3233.170 ;
        RECT 2686.630 3053.590 2687.810 3054.770 ;
        RECT 2688.230 3053.590 2689.410 3054.770 ;
        RECT 2686.630 3051.990 2687.810 3053.170 ;
        RECT 2688.230 3051.990 2689.410 3053.170 ;
        RECT 2686.630 2873.590 2687.810 2874.770 ;
        RECT 2688.230 2873.590 2689.410 2874.770 ;
        RECT 2686.630 2871.990 2687.810 2873.170 ;
        RECT 2688.230 2871.990 2689.410 2873.170 ;
        RECT 2686.630 2693.590 2687.810 2694.770 ;
        RECT 2688.230 2693.590 2689.410 2694.770 ;
        RECT 2686.630 2691.990 2687.810 2693.170 ;
        RECT 2688.230 2691.990 2689.410 2693.170 ;
        RECT 2686.630 2513.590 2687.810 2514.770 ;
        RECT 2688.230 2513.590 2689.410 2514.770 ;
        RECT 2686.630 2511.990 2687.810 2513.170 ;
        RECT 2688.230 2511.990 2689.410 2513.170 ;
        RECT 2686.630 2333.590 2687.810 2334.770 ;
        RECT 2688.230 2333.590 2689.410 2334.770 ;
        RECT 2686.630 2331.990 2687.810 2333.170 ;
        RECT 2688.230 2331.990 2689.410 2333.170 ;
        RECT 2686.630 2153.590 2687.810 2154.770 ;
        RECT 2688.230 2153.590 2689.410 2154.770 ;
        RECT 2686.630 2151.990 2687.810 2153.170 ;
        RECT 2688.230 2151.990 2689.410 2153.170 ;
        RECT 2686.630 1973.590 2687.810 1974.770 ;
        RECT 2688.230 1973.590 2689.410 1974.770 ;
        RECT 2686.630 1971.990 2687.810 1973.170 ;
        RECT 2688.230 1971.990 2689.410 1973.170 ;
        RECT 2686.630 1793.590 2687.810 1794.770 ;
        RECT 2688.230 1793.590 2689.410 1794.770 ;
        RECT 2686.630 1791.990 2687.810 1793.170 ;
        RECT 2688.230 1791.990 2689.410 1793.170 ;
        RECT 2686.630 1613.590 2687.810 1614.770 ;
        RECT 2688.230 1613.590 2689.410 1614.770 ;
        RECT 2686.630 1611.990 2687.810 1613.170 ;
        RECT 2688.230 1611.990 2689.410 1613.170 ;
        RECT 2686.630 1433.590 2687.810 1434.770 ;
        RECT 2688.230 1433.590 2689.410 1434.770 ;
        RECT 2686.630 1431.990 2687.810 1433.170 ;
        RECT 2688.230 1431.990 2689.410 1433.170 ;
        RECT 2686.630 1253.590 2687.810 1254.770 ;
        RECT 2688.230 1253.590 2689.410 1254.770 ;
        RECT 2686.630 1251.990 2687.810 1253.170 ;
        RECT 2688.230 1251.990 2689.410 1253.170 ;
        RECT 2686.630 1073.590 2687.810 1074.770 ;
        RECT 2688.230 1073.590 2689.410 1074.770 ;
        RECT 2686.630 1071.990 2687.810 1073.170 ;
        RECT 2688.230 1071.990 2689.410 1073.170 ;
        RECT 2686.630 893.590 2687.810 894.770 ;
        RECT 2688.230 893.590 2689.410 894.770 ;
        RECT 2686.630 891.990 2687.810 893.170 ;
        RECT 2688.230 891.990 2689.410 893.170 ;
        RECT 2686.630 713.590 2687.810 714.770 ;
        RECT 2688.230 713.590 2689.410 714.770 ;
        RECT 2686.630 711.990 2687.810 713.170 ;
        RECT 2688.230 711.990 2689.410 713.170 ;
        RECT 2686.630 533.590 2687.810 534.770 ;
        RECT 2688.230 533.590 2689.410 534.770 ;
        RECT 2686.630 531.990 2687.810 533.170 ;
        RECT 2688.230 531.990 2689.410 533.170 ;
        RECT 2686.630 353.590 2687.810 354.770 ;
        RECT 2688.230 353.590 2689.410 354.770 ;
        RECT 2686.630 351.990 2687.810 353.170 ;
        RECT 2688.230 351.990 2689.410 353.170 ;
        RECT 2686.630 173.590 2687.810 174.770 ;
        RECT 2688.230 173.590 2689.410 174.770 ;
        RECT 2686.630 171.990 2687.810 173.170 ;
        RECT 2688.230 171.990 2689.410 173.170 ;
        RECT 2686.630 -36.510 2687.810 -35.330 ;
        RECT 2688.230 -36.510 2689.410 -35.330 ;
        RECT 2686.630 -38.110 2687.810 -36.930 ;
        RECT 2688.230 -38.110 2689.410 -36.930 ;
        RECT 2866.630 3556.610 2867.810 3557.790 ;
        RECT 2868.230 3556.610 2869.410 3557.790 ;
        RECT 2866.630 3555.010 2867.810 3556.190 ;
        RECT 2868.230 3555.010 2869.410 3556.190 ;
        RECT 2866.630 3413.590 2867.810 3414.770 ;
        RECT 2868.230 3413.590 2869.410 3414.770 ;
        RECT 2866.630 3411.990 2867.810 3413.170 ;
        RECT 2868.230 3411.990 2869.410 3413.170 ;
        RECT 2866.630 3233.590 2867.810 3234.770 ;
        RECT 2868.230 3233.590 2869.410 3234.770 ;
        RECT 2866.630 3231.990 2867.810 3233.170 ;
        RECT 2868.230 3231.990 2869.410 3233.170 ;
        RECT 2866.630 3053.590 2867.810 3054.770 ;
        RECT 2868.230 3053.590 2869.410 3054.770 ;
        RECT 2866.630 3051.990 2867.810 3053.170 ;
        RECT 2868.230 3051.990 2869.410 3053.170 ;
        RECT 2866.630 2873.590 2867.810 2874.770 ;
        RECT 2868.230 2873.590 2869.410 2874.770 ;
        RECT 2866.630 2871.990 2867.810 2873.170 ;
        RECT 2868.230 2871.990 2869.410 2873.170 ;
        RECT 2866.630 2693.590 2867.810 2694.770 ;
        RECT 2868.230 2693.590 2869.410 2694.770 ;
        RECT 2866.630 2691.990 2867.810 2693.170 ;
        RECT 2868.230 2691.990 2869.410 2693.170 ;
        RECT 2866.630 2513.590 2867.810 2514.770 ;
        RECT 2868.230 2513.590 2869.410 2514.770 ;
        RECT 2866.630 2511.990 2867.810 2513.170 ;
        RECT 2868.230 2511.990 2869.410 2513.170 ;
        RECT 2866.630 2333.590 2867.810 2334.770 ;
        RECT 2868.230 2333.590 2869.410 2334.770 ;
        RECT 2866.630 2331.990 2867.810 2333.170 ;
        RECT 2868.230 2331.990 2869.410 2333.170 ;
        RECT 2866.630 2153.590 2867.810 2154.770 ;
        RECT 2868.230 2153.590 2869.410 2154.770 ;
        RECT 2866.630 2151.990 2867.810 2153.170 ;
        RECT 2868.230 2151.990 2869.410 2153.170 ;
        RECT 2866.630 1973.590 2867.810 1974.770 ;
        RECT 2868.230 1973.590 2869.410 1974.770 ;
        RECT 2866.630 1971.990 2867.810 1973.170 ;
        RECT 2868.230 1971.990 2869.410 1973.170 ;
        RECT 2866.630 1793.590 2867.810 1794.770 ;
        RECT 2868.230 1793.590 2869.410 1794.770 ;
        RECT 2866.630 1791.990 2867.810 1793.170 ;
        RECT 2868.230 1791.990 2869.410 1793.170 ;
        RECT 2866.630 1613.590 2867.810 1614.770 ;
        RECT 2868.230 1613.590 2869.410 1614.770 ;
        RECT 2866.630 1611.990 2867.810 1613.170 ;
        RECT 2868.230 1611.990 2869.410 1613.170 ;
        RECT 2866.630 1433.590 2867.810 1434.770 ;
        RECT 2868.230 1433.590 2869.410 1434.770 ;
        RECT 2866.630 1431.990 2867.810 1433.170 ;
        RECT 2868.230 1431.990 2869.410 1433.170 ;
        RECT 2866.630 1253.590 2867.810 1254.770 ;
        RECT 2868.230 1253.590 2869.410 1254.770 ;
        RECT 2866.630 1251.990 2867.810 1253.170 ;
        RECT 2868.230 1251.990 2869.410 1253.170 ;
        RECT 2866.630 1073.590 2867.810 1074.770 ;
        RECT 2868.230 1073.590 2869.410 1074.770 ;
        RECT 2866.630 1071.990 2867.810 1073.170 ;
        RECT 2868.230 1071.990 2869.410 1073.170 ;
        RECT 2866.630 893.590 2867.810 894.770 ;
        RECT 2868.230 893.590 2869.410 894.770 ;
        RECT 2866.630 891.990 2867.810 893.170 ;
        RECT 2868.230 891.990 2869.410 893.170 ;
        RECT 2866.630 713.590 2867.810 714.770 ;
        RECT 2868.230 713.590 2869.410 714.770 ;
        RECT 2866.630 711.990 2867.810 713.170 ;
        RECT 2868.230 711.990 2869.410 713.170 ;
        RECT 2866.630 533.590 2867.810 534.770 ;
        RECT 2868.230 533.590 2869.410 534.770 ;
        RECT 2866.630 531.990 2867.810 533.170 ;
        RECT 2868.230 531.990 2869.410 533.170 ;
        RECT 2866.630 353.590 2867.810 354.770 ;
        RECT 2868.230 353.590 2869.410 354.770 ;
        RECT 2866.630 351.990 2867.810 353.170 ;
        RECT 2868.230 351.990 2869.410 353.170 ;
        RECT 2866.630 173.590 2867.810 174.770 ;
        RECT 2868.230 173.590 2869.410 174.770 ;
        RECT 2866.630 171.990 2867.810 173.170 ;
        RECT 2868.230 171.990 2869.410 173.170 ;
        RECT 2866.630 -36.510 2867.810 -35.330 ;
        RECT 2868.230 -36.510 2869.410 -35.330 ;
        RECT 2866.630 -38.110 2867.810 -36.930 ;
        RECT 2868.230 -38.110 2869.410 -36.930 ;
        RECT 2960.310 3556.610 2961.490 3557.790 ;
        RECT 2961.910 3556.610 2963.090 3557.790 ;
        RECT 2960.310 3555.010 2961.490 3556.190 ;
        RECT 2961.910 3555.010 2963.090 3556.190 ;
        RECT 2960.310 3413.590 2961.490 3414.770 ;
        RECT 2961.910 3413.590 2963.090 3414.770 ;
        RECT 2960.310 3411.990 2961.490 3413.170 ;
        RECT 2961.910 3411.990 2963.090 3413.170 ;
        RECT 2960.310 3233.590 2961.490 3234.770 ;
        RECT 2961.910 3233.590 2963.090 3234.770 ;
        RECT 2960.310 3231.990 2961.490 3233.170 ;
        RECT 2961.910 3231.990 2963.090 3233.170 ;
        RECT 2960.310 3053.590 2961.490 3054.770 ;
        RECT 2961.910 3053.590 2963.090 3054.770 ;
        RECT 2960.310 3051.990 2961.490 3053.170 ;
        RECT 2961.910 3051.990 2963.090 3053.170 ;
        RECT 2960.310 2873.590 2961.490 2874.770 ;
        RECT 2961.910 2873.590 2963.090 2874.770 ;
        RECT 2960.310 2871.990 2961.490 2873.170 ;
        RECT 2961.910 2871.990 2963.090 2873.170 ;
        RECT 2960.310 2693.590 2961.490 2694.770 ;
        RECT 2961.910 2693.590 2963.090 2694.770 ;
        RECT 2960.310 2691.990 2961.490 2693.170 ;
        RECT 2961.910 2691.990 2963.090 2693.170 ;
        RECT 2960.310 2513.590 2961.490 2514.770 ;
        RECT 2961.910 2513.590 2963.090 2514.770 ;
        RECT 2960.310 2511.990 2961.490 2513.170 ;
        RECT 2961.910 2511.990 2963.090 2513.170 ;
        RECT 2960.310 2333.590 2961.490 2334.770 ;
        RECT 2961.910 2333.590 2963.090 2334.770 ;
        RECT 2960.310 2331.990 2961.490 2333.170 ;
        RECT 2961.910 2331.990 2963.090 2333.170 ;
        RECT 2960.310 2153.590 2961.490 2154.770 ;
        RECT 2961.910 2153.590 2963.090 2154.770 ;
        RECT 2960.310 2151.990 2961.490 2153.170 ;
        RECT 2961.910 2151.990 2963.090 2153.170 ;
        RECT 2960.310 1973.590 2961.490 1974.770 ;
        RECT 2961.910 1973.590 2963.090 1974.770 ;
        RECT 2960.310 1971.990 2961.490 1973.170 ;
        RECT 2961.910 1971.990 2963.090 1973.170 ;
        RECT 2960.310 1793.590 2961.490 1794.770 ;
        RECT 2961.910 1793.590 2963.090 1794.770 ;
        RECT 2960.310 1791.990 2961.490 1793.170 ;
        RECT 2961.910 1791.990 2963.090 1793.170 ;
        RECT 2960.310 1613.590 2961.490 1614.770 ;
        RECT 2961.910 1613.590 2963.090 1614.770 ;
        RECT 2960.310 1611.990 2961.490 1613.170 ;
        RECT 2961.910 1611.990 2963.090 1613.170 ;
        RECT 2960.310 1433.590 2961.490 1434.770 ;
        RECT 2961.910 1433.590 2963.090 1434.770 ;
        RECT 2960.310 1431.990 2961.490 1433.170 ;
        RECT 2961.910 1431.990 2963.090 1433.170 ;
        RECT 2960.310 1253.590 2961.490 1254.770 ;
        RECT 2961.910 1253.590 2963.090 1254.770 ;
        RECT 2960.310 1251.990 2961.490 1253.170 ;
        RECT 2961.910 1251.990 2963.090 1253.170 ;
        RECT 2960.310 1073.590 2961.490 1074.770 ;
        RECT 2961.910 1073.590 2963.090 1074.770 ;
        RECT 2960.310 1071.990 2961.490 1073.170 ;
        RECT 2961.910 1071.990 2963.090 1073.170 ;
        RECT 2960.310 893.590 2961.490 894.770 ;
        RECT 2961.910 893.590 2963.090 894.770 ;
        RECT 2960.310 891.990 2961.490 893.170 ;
        RECT 2961.910 891.990 2963.090 893.170 ;
        RECT 2960.310 713.590 2961.490 714.770 ;
        RECT 2961.910 713.590 2963.090 714.770 ;
        RECT 2960.310 711.990 2961.490 713.170 ;
        RECT 2961.910 711.990 2963.090 713.170 ;
        RECT 2960.310 533.590 2961.490 534.770 ;
        RECT 2961.910 533.590 2963.090 534.770 ;
        RECT 2960.310 531.990 2961.490 533.170 ;
        RECT 2961.910 531.990 2963.090 533.170 ;
        RECT 2960.310 353.590 2961.490 354.770 ;
        RECT 2961.910 353.590 2963.090 354.770 ;
        RECT 2960.310 351.990 2961.490 353.170 ;
        RECT 2961.910 351.990 2963.090 353.170 ;
        RECT 2960.310 173.590 2961.490 174.770 ;
        RECT 2961.910 173.590 2963.090 174.770 ;
        RECT 2960.310 171.990 2961.490 173.170 ;
        RECT 2961.910 171.990 2963.090 173.170 ;
        RECT 2960.310 -36.510 2961.490 -35.330 ;
        RECT 2961.910 -36.510 2963.090 -35.330 ;
        RECT 2960.310 -38.110 2961.490 -36.930 ;
        RECT 2961.910 -38.110 2963.090 -36.930 ;
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
        RECT -43.630 3411.830 2963.250 3414.930 ;
        RECT -43.630 3231.830 2963.250 3234.930 ;
        RECT -43.630 3051.830 2963.250 3054.930 ;
        RECT -43.630 2871.830 2963.250 2874.930 ;
        RECT -43.630 2691.830 2963.250 2694.930 ;
        RECT -43.630 2511.830 2963.250 2514.930 ;
        RECT -43.630 2331.830 2963.250 2334.930 ;
        RECT -43.630 2151.830 2963.250 2154.930 ;
        RECT -43.630 1971.830 2963.250 1974.930 ;
        RECT -43.630 1791.830 2963.250 1794.930 ;
        RECT -43.630 1611.830 2963.250 1614.930 ;
        RECT -43.630 1431.830 2963.250 1434.930 ;
        RECT -43.630 1251.830 2963.250 1254.930 ;
        RECT -43.630 1071.830 2963.250 1074.930 ;
        RECT -43.630 891.830 2963.250 894.930 ;
        RECT -43.630 711.830 2963.250 714.930 ;
        RECT -43.630 531.830 2963.250 534.930 ;
        RECT -43.630 351.830 2963.250 354.930 ;
        RECT -43.630 171.830 2963.250 174.930 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
        RECT 31.470 -38.270 34.570 3557.950 ;
        RECT 211.470 -38.270 214.570 3557.950 ;
        RECT 391.470 810.000 394.570 3557.950 ;
        RECT 571.470 810.000 574.570 3557.950 ;
        RECT 497.840 510.640 499.440 788.560 ;
        RECT 651.440 510.640 653.040 788.560 ;
        RECT 391.470 -38.270 394.570 490.000 ;
        RECT 571.470 -38.270 574.570 490.000 ;
        RECT 751.470 -38.270 754.570 3557.950 ;
        RECT 931.470 -38.270 934.570 3557.950 ;
        RECT 1111.470 -38.270 1114.570 3557.950 ;
        RECT 1291.470 -38.270 1294.570 3557.950 ;
        RECT 1471.470 -38.270 1474.570 3557.950 ;
        RECT 1651.470 -38.270 1654.570 3557.950 ;
        RECT 1831.470 -38.270 1834.570 3557.950 ;
        RECT 2011.470 -38.270 2014.570 3557.950 ;
        RECT 2191.470 -38.270 2194.570 3557.950 ;
        RECT 2371.470 -38.270 2374.570 3557.950 ;
        RECT 2551.470 -38.270 2554.570 3557.950 ;
        RECT 2731.470 -38.270 2734.570 3557.950 ;
        RECT 2911.470 -38.270 2914.570 3557.950 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
      LAYER via4 ;
        RECT -14.670 3527.810 -13.490 3528.990 ;
        RECT -13.070 3527.810 -11.890 3528.990 ;
        RECT -14.670 3526.210 -13.490 3527.390 ;
        RECT -13.070 3526.210 -11.890 3527.390 ;
        RECT -14.670 3458.590 -13.490 3459.770 ;
        RECT -13.070 3458.590 -11.890 3459.770 ;
        RECT -14.670 3456.990 -13.490 3458.170 ;
        RECT -13.070 3456.990 -11.890 3458.170 ;
        RECT -14.670 3278.590 -13.490 3279.770 ;
        RECT -13.070 3278.590 -11.890 3279.770 ;
        RECT -14.670 3276.990 -13.490 3278.170 ;
        RECT -13.070 3276.990 -11.890 3278.170 ;
        RECT -14.670 3098.590 -13.490 3099.770 ;
        RECT -13.070 3098.590 -11.890 3099.770 ;
        RECT -14.670 3096.990 -13.490 3098.170 ;
        RECT -13.070 3096.990 -11.890 3098.170 ;
        RECT -14.670 2918.590 -13.490 2919.770 ;
        RECT -13.070 2918.590 -11.890 2919.770 ;
        RECT -14.670 2916.990 -13.490 2918.170 ;
        RECT -13.070 2916.990 -11.890 2918.170 ;
        RECT -14.670 2738.590 -13.490 2739.770 ;
        RECT -13.070 2738.590 -11.890 2739.770 ;
        RECT -14.670 2736.990 -13.490 2738.170 ;
        RECT -13.070 2736.990 -11.890 2738.170 ;
        RECT -14.670 2558.590 -13.490 2559.770 ;
        RECT -13.070 2558.590 -11.890 2559.770 ;
        RECT -14.670 2556.990 -13.490 2558.170 ;
        RECT -13.070 2556.990 -11.890 2558.170 ;
        RECT -14.670 2378.590 -13.490 2379.770 ;
        RECT -13.070 2378.590 -11.890 2379.770 ;
        RECT -14.670 2376.990 -13.490 2378.170 ;
        RECT -13.070 2376.990 -11.890 2378.170 ;
        RECT -14.670 2198.590 -13.490 2199.770 ;
        RECT -13.070 2198.590 -11.890 2199.770 ;
        RECT -14.670 2196.990 -13.490 2198.170 ;
        RECT -13.070 2196.990 -11.890 2198.170 ;
        RECT -14.670 2018.590 -13.490 2019.770 ;
        RECT -13.070 2018.590 -11.890 2019.770 ;
        RECT -14.670 2016.990 -13.490 2018.170 ;
        RECT -13.070 2016.990 -11.890 2018.170 ;
        RECT -14.670 1838.590 -13.490 1839.770 ;
        RECT -13.070 1838.590 -11.890 1839.770 ;
        RECT -14.670 1836.990 -13.490 1838.170 ;
        RECT -13.070 1836.990 -11.890 1838.170 ;
        RECT -14.670 1658.590 -13.490 1659.770 ;
        RECT -13.070 1658.590 -11.890 1659.770 ;
        RECT -14.670 1656.990 -13.490 1658.170 ;
        RECT -13.070 1656.990 -11.890 1658.170 ;
        RECT -14.670 1478.590 -13.490 1479.770 ;
        RECT -13.070 1478.590 -11.890 1479.770 ;
        RECT -14.670 1476.990 -13.490 1478.170 ;
        RECT -13.070 1476.990 -11.890 1478.170 ;
        RECT -14.670 1298.590 -13.490 1299.770 ;
        RECT -13.070 1298.590 -11.890 1299.770 ;
        RECT -14.670 1296.990 -13.490 1298.170 ;
        RECT -13.070 1296.990 -11.890 1298.170 ;
        RECT -14.670 1118.590 -13.490 1119.770 ;
        RECT -13.070 1118.590 -11.890 1119.770 ;
        RECT -14.670 1116.990 -13.490 1118.170 ;
        RECT -13.070 1116.990 -11.890 1118.170 ;
        RECT -14.670 938.590 -13.490 939.770 ;
        RECT -13.070 938.590 -11.890 939.770 ;
        RECT -14.670 936.990 -13.490 938.170 ;
        RECT -13.070 936.990 -11.890 938.170 ;
        RECT -14.670 758.590 -13.490 759.770 ;
        RECT -13.070 758.590 -11.890 759.770 ;
        RECT -14.670 756.990 -13.490 758.170 ;
        RECT -13.070 756.990 -11.890 758.170 ;
        RECT -14.670 578.590 -13.490 579.770 ;
        RECT -13.070 578.590 -11.890 579.770 ;
        RECT -14.670 576.990 -13.490 578.170 ;
        RECT -13.070 576.990 -11.890 578.170 ;
        RECT -14.670 398.590 -13.490 399.770 ;
        RECT -13.070 398.590 -11.890 399.770 ;
        RECT -14.670 396.990 -13.490 398.170 ;
        RECT -13.070 396.990 -11.890 398.170 ;
        RECT -14.670 218.590 -13.490 219.770 ;
        RECT -13.070 218.590 -11.890 219.770 ;
        RECT -14.670 216.990 -13.490 218.170 ;
        RECT -13.070 216.990 -11.890 218.170 ;
        RECT -14.670 38.590 -13.490 39.770 ;
        RECT -13.070 38.590 -11.890 39.770 ;
        RECT -14.670 36.990 -13.490 38.170 ;
        RECT -13.070 36.990 -11.890 38.170 ;
        RECT -14.670 -7.710 -13.490 -6.530 ;
        RECT -13.070 -7.710 -11.890 -6.530 ;
        RECT -14.670 -9.310 -13.490 -8.130 ;
        RECT -13.070 -9.310 -11.890 -8.130 ;
        RECT 31.630 3527.810 32.810 3528.990 ;
        RECT 33.230 3527.810 34.410 3528.990 ;
        RECT 31.630 3526.210 32.810 3527.390 ;
        RECT 33.230 3526.210 34.410 3527.390 ;
        RECT 31.630 3458.590 32.810 3459.770 ;
        RECT 33.230 3458.590 34.410 3459.770 ;
        RECT 31.630 3456.990 32.810 3458.170 ;
        RECT 33.230 3456.990 34.410 3458.170 ;
        RECT 31.630 3278.590 32.810 3279.770 ;
        RECT 33.230 3278.590 34.410 3279.770 ;
        RECT 31.630 3276.990 32.810 3278.170 ;
        RECT 33.230 3276.990 34.410 3278.170 ;
        RECT 31.630 3098.590 32.810 3099.770 ;
        RECT 33.230 3098.590 34.410 3099.770 ;
        RECT 31.630 3096.990 32.810 3098.170 ;
        RECT 33.230 3096.990 34.410 3098.170 ;
        RECT 31.630 2918.590 32.810 2919.770 ;
        RECT 33.230 2918.590 34.410 2919.770 ;
        RECT 31.630 2916.990 32.810 2918.170 ;
        RECT 33.230 2916.990 34.410 2918.170 ;
        RECT 31.630 2738.590 32.810 2739.770 ;
        RECT 33.230 2738.590 34.410 2739.770 ;
        RECT 31.630 2736.990 32.810 2738.170 ;
        RECT 33.230 2736.990 34.410 2738.170 ;
        RECT 31.630 2558.590 32.810 2559.770 ;
        RECT 33.230 2558.590 34.410 2559.770 ;
        RECT 31.630 2556.990 32.810 2558.170 ;
        RECT 33.230 2556.990 34.410 2558.170 ;
        RECT 31.630 2378.590 32.810 2379.770 ;
        RECT 33.230 2378.590 34.410 2379.770 ;
        RECT 31.630 2376.990 32.810 2378.170 ;
        RECT 33.230 2376.990 34.410 2378.170 ;
        RECT 31.630 2198.590 32.810 2199.770 ;
        RECT 33.230 2198.590 34.410 2199.770 ;
        RECT 31.630 2196.990 32.810 2198.170 ;
        RECT 33.230 2196.990 34.410 2198.170 ;
        RECT 31.630 2018.590 32.810 2019.770 ;
        RECT 33.230 2018.590 34.410 2019.770 ;
        RECT 31.630 2016.990 32.810 2018.170 ;
        RECT 33.230 2016.990 34.410 2018.170 ;
        RECT 31.630 1838.590 32.810 1839.770 ;
        RECT 33.230 1838.590 34.410 1839.770 ;
        RECT 31.630 1836.990 32.810 1838.170 ;
        RECT 33.230 1836.990 34.410 1838.170 ;
        RECT 31.630 1658.590 32.810 1659.770 ;
        RECT 33.230 1658.590 34.410 1659.770 ;
        RECT 31.630 1656.990 32.810 1658.170 ;
        RECT 33.230 1656.990 34.410 1658.170 ;
        RECT 31.630 1478.590 32.810 1479.770 ;
        RECT 33.230 1478.590 34.410 1479.770 ;
        RECT 31.630 1476.990 32.810 1478.170 ;
        RECT 33.230 1476.990 34.410 1478.170 ;
        RECT 31.630 1298.590 32.810 1299.770 ;
        RECT 33.230 1298.590 34.410 1299.770 ;
        RECT 31.630 1296.990 32.810 1298.170 ;
        RECT 33.230 1296.990 34.410 1298.170 ;
        RECT 31.630 1118.590 32.810 1119.770 ;
        RECT 33.230 1118.590 34.410 1119.770 ;
        RECT 31.630 1116.990 32.810 1118.170 ;
        RECT 33.230 1116.990 34.410 1118.170 ;
        RECT 31.630 938.590 32.810 939.770 ;
        RECT 33.230 938.590 34.410 939.770 ;
        RECT 31.630 936.990 32.810 938.170 ;
        RECT 33.230 936.990 34.410 938.170 ;
        RECT 31.630 758.590 32.810 759.770 ;
        RECT 33.230 758.590 34.410 759.770 ;
        RECT 31.630 756.990 32.810 758.170 ;
        RECT 33.230 756.990 34.410 758.170 ;
        RECT 31.630 578.590 32.810 579.770 ;
        RECT 33.230 578.590 34.410 579.770 ;
        RECT 31.630 576.990 32.810 578.170 ;
        RECT 33.230 576.990 34.410 578.170 ;
        RECT 31.630 398.590 32.810 399.770 ;
        RECT 33.230 398.590 34.410 399.770 ;
        RECT 31.630 396.990 32.810 398.170 ;
        RECT 33.230 396.990 34.410 398.170 ;
        RECT 31.630 218.590 32.810 219.770 ;
        RECT 33.230 218.590 34.410 219.770 ;
        RECT 31.630 216.990 32.810 218.170 ;
        RECT 33.230 216.990 34.410 218.170 ;
        RECT 31.630 38.590 32.810 39.770 ;
        RECT 33.230 38.590 34.410 39.770 ;
        RECT 31.630 36.990 32.810 38.170 ;
        RECT 33.230 36.990 34.410 38.170 ;
        RECT 31.630 -7.710 32.810 -6.530 ;
        RECT 33.230 -7.710 34.410 -6.530 ;
        RECT 31.630 -9.310 32.810 -8.130 ;
        RECT 33.230 -9.310 34.410 -8.130 ;
        RECT 211.630 3527.810 212.810 3528.990 ;
        RECT 213.230 3527.810 214.410 3528.990 ;
        RECT 211.630 3526.210 212.810 3527.390 ;
        RECT 213.230 3526.210 214.410 3527.390 ;
        RECT 211.630 3458.590 212.810 3459.770 ;
        RECT 213.230 3458.590 214.410 3459.770 ;
        RECT 211.630 3456.990 212.810 3458.170 ;
        RECT 213.230 3456.990 214.410 3458.170 ;
        RECT 211.630 3278.590 212.810 3279.770 ;
        RECT 213.230 3278.590 214.410 3279.770 ;
        RECT 211.630 3276.990 212.810 3278.170 ;
        RECT 213.230 3276.990 214.410 3278.170 ;
        RECT 211.630 3098.590 212.810 3099.770 ;
        RECT 213.230 3098.590 214.410 3099.770 ;
        RECT 211.630 3096.990 212.810 3098.170 ;
        RECT 213.230 3096.990 214.410 3098.170 ;
        RECT 211.630 2918.590 212.810 2919.770 ;
        RECT 213.230 2918.590 214.410 2919.770 ;
        RECT 211.630 2916.990 212.810 2918.170 ;
        RECT 213.230 2916.990 214.410 2918.170 ;
        RECT 211.630 2738.590 212.810 2739.770 ;
        RECT 213.230 2738.590 214.410 2739.770 ;
        RECT 211.630 2736.990 212.810 2738.170 ;
        RECT 213.230 2736.990 214.410 2738.170 ;
        RECT 211.630 2558.590 212.810 2559.770 ;
        RECT 213.230 2558.590 214.410 2559.770 ;
        RECT 211.630 2556.990 212.810 2558.170 ;
        RECT 213.230 2556.990 214.410 2558.170 ;
        RECT 211.630 2378.590 212.810 2379.770 ;
        RECT 213.230 2378.590 214.410 2379.770 ;
        RECT 211.630 2376.990 212.810 2378.170 ;
        RECT 213.230 2376.990 214.410 2378.170 ;
        RECT 211.630 2198.590 212.810 2199.770 ;
        RECT 213.230 2198.590 214.410 2199.770 ;
        RECT 211.630 2196.990 212.810 2198.170 ;
        RECT 213.230 2196.990 214.410 2198.170 ;
        RECT 211.630 2018.590 212.810 2019.770 ;
        RECT 213.230 2018.590 214.410 2019.770 ;
        RECT 211.630 2016.990 212.810 2018.170 ;
        RECT 213.230 2016.990 214.410 2018.170 ;
        RECT 211.630 1838.590 212.810 1839.770 ;
        RECT 213.230 1838.590 214.410 1839.770 ;
        RECT 211.630 1836.990 212.810 1838.170 ;
        RECT 213.230 1836.990 214.410 1838.170 ;
        RECT 211.630 1658.590 212.810 1659.770 ;
        RECT 213.230 1658.590 214.410 1659.770 ;
        RECT 211.630 1656.990 212.810 1658.170 ;
        RECT 213.230 1656.990 214.410 1658.170 ;
        RECT 211.630 1478.590 212.810 1479.770 ;
        RECT 213.230 1478.590 214.410 1479.770 ;
        RECT 211.630 1476.990 212.810 1478.170 ;
        RECT 213.230 1476.990 214.410 1478.170 ;
        RECT 211.630 1298.590 212.810 1299.770 ;
        RECT 213.230 1298.590 214.410 1299.770 ;
        RECT 211.630 1296.990 212.810 1298.170 ;
        RECT 213.230 1296.990 214.410 1298.170 ;
        RECT 211.630 1118.590 212.810 1119.770 ;
        RECT 213.230 1118.590 214.410 1119.770 ;
        RECT 211.630 1116.990 212.810 1118.170 ;
        RECT 213.230 1116.990 214.410 1118.170 ;
        RECT 211.630 938.590 212.810 939.770 ;
        RECT 213.230 938.590 214.410 939.770 ;
        RECT 211.630 936.990 212.810 938.170 ;
        RECT 213.230 936.990 214.410 938.170 ;
        RECT 391.630 3527.810 392.810 3528.990 ;
        RECT 393.230 3527.810 394.410 3528.990 ;
        RECT 391.630 3526.210 392.810 3527.390 ;
        RECT 393.230 3526.210 394.410 3527.390 ;
        RECT 391.630 3458.590 392.810 3459.770 ;
        RECT 393.230 3458.590 394.410 3459.770 ;
        RECT 391.630 3456.990 392.810 3458.170 ;
        RECT 393.230 3456.990 394.410 3458.170 ;
        RECT 391.630 3278.590 392.810 3279.770 ;
        RECT 393.230 3278.590 394.410 3279.770 ;
        RECT 391.630 3276.990 392.810 3278.170 ;
        RECT 393.230 3276.990 394.410 3278.170 ;
        RECT 391.630 3098.590 392.810 3099.770 ;
        RECT 393.230 3098.590 394.410 3099.770 ;
        RECT 391.630 3096.990 392.810 3098.170 ;
        RECT 393.230 3096.990 394.410 3098.170 ;
        RECT 391.630 2918.590 392.810 2919.770 ;
        RECT 393.230 2918.590 394.410 2919.770 ;
        RECT 391.630 2916.990 392.810 2918.170 ;
        RECT 393.230 2916.990 394.410 2918.170 ;
        RECT 391.630 2738.590 392.810 2739.770 ;
        RECT 393.230 2738.590 394.410 2739.770 ;
        RECT 391.630 2736.990 392.810 2738.170 ;
        RECT 393.230 2736.990 394.410 2738.170 ;
        RECT 391.630 2558.590 392.810 2559.770 ;
        RECT 393.230 2558.590 394.410 2559.770 ;
        RECT 391.630 2556.990 392.810 2558.170 ;
        RECT 393.230 2556.990 394.410 2558.170 ;
        RECT 391.630 2378.590 392.810 2379.770 ;
        RECT 393.230 2378.590 394.410 2379.770 ;
        RECT 391.630 2376.990 392.810 2378.170 ;
        RECT 393.230 2376.990 394.410 2378.170 ;
        RECT 391.630 2198.590 392.810 2199.770 ;
        RECT 393.230 2198.590 394.410 2199.770 ;
        RECT 391.630 2196.990 392.810 2198.170 ;
        RECT 393.230 2196.990 394.410 2198.170 ;
        RECT 391.630 2018.590 392.810 2019.770 ;
        RECT 393.230 2018.590 394.410 2019.770 ;
        RECT 391.630 2016.990 392.810 2018.170 ;
        RECT 393.230 2016.990 394.410 2018.170 ;
        RECT 391.630 1838.590 392.810 1839.770 ;
        RECT 393.230 1838.590 394.410 1839.770 ;
        RECT 391.630 1836.990 392.810 1838.170 ;
        RECT 393.230 1836.990 394.410 1838.170 ;
        RECT 391.630 1658.590 392.810 1659.770 ;
        RECT 393.230 1658.590 394.410 1659.770 ;
        RECT 391.630 1656.990 392.810 1658.170 ;
        RECT 393.230 1656.990 394.410 1658.170 ;
        RECT 391.630 1478.590 392.810 1479.770 ;
        RECT 393.230 1478.590 394.410 1479.770 ;
        RECT 391.630 1476.990 392.810 1478.170 ;
        RECT 393.230 1476.990 394.410 1478.170 ;
        RECT 391.630 1298.590 392.810 1299.770 ;
        RECT 393.230 1298.590 394.410 1299.770 ;
        RECT 391.630 1296.990 392.810 1298.170 ;
        RECT 393.230 1296.990 394.410 1298.170 ;
        RECT 391.630 1118.590 392.810 1119.770 ;
        RECT 393.230 1118.590 394.410 1119.770 ;
        RECT 391.630 1116.990 392.810 1118.170 ;
        RECT 393.230 1116.990 394.410 1118.170 ;
        RECT 391.630 938.590 392.810 939.770 ;
        RECT 393.230 938.590 394.410 939.770 ;
        RECT 391.630 936.990 392.810 938.170 ;
        RECT 393.230 936.990 394.410 938.170 ;
        RECT 571.630 3527.810 572.810 3528.990 ;
        RECT 573.230 3527.810 574.410 3528.990 ;
        RECT 571.630 3526.210 572.810 3527.390 ;
        RECT 573.230 3526.210 574.410 3527.390 ;
        RECT 571.630 3458.590 572.810 3459.770 ;
        RECT 573.230 3458.590 574.410 3459.770 ;
        RECT 571.630 3456.990 572.810 3458.170 ;
        RECT 573.230 3456.990 574.410 3458.170 ;
        RECT 571.630 3278.590 572.810 3279.770 ;
        RECT 573.230 3278.590 574.410 3279.770 ;
        RECT 571.630 3276.990 572.810 3278.170 ;
        RECT 573.230 3276.990 574.410 3278.170 ;
        RECT 571.630 3098.590 572.810 3099.770 ;
        RECT 573.230 3098.590 574.410 3099.770 ;
        RECT 571.630 3096.990 572.810 3098.170 ;
        RECT 573.230 3096.990 574.410 3098.170 ;
        RECT 571.630 2918.590 572.810 2919.770 ;
        RECT 573.230 2918.590 574.410 2919.770 ;
        RECT 571.630 2916.990 572.810 2918.170 ;
        RECT 573.230 2916.990 574.410 2918.170 ;
        RECT 571.630 2738.590 572.810 2739.770 ;
        RECT 573.230 2738.590 574.410 2739.770 ;
        RECT 571.630 2736.990 572.810 2738.170 ;
        RECT 573.230 2736.990 574.410 2738.170 ;
        RECT 571.630 2558.590 572.810 2559.770 ;
        RECT 573.230 2558.590 574.410 2559.770 ;
        RECT 571.630 2556.990 572.810 2558.170 ;
        RECT 573.230 2556.990 574.410 2558.170 ;
        RECT 571.630 2378.590 572.810 2379.770 ;
        RECT 573.230 2378.590 574.410 2379.770 ;
        RECT 571.630 2376.990 572.810 2378.170 ;
        RECT 573.230 2376.990 574.410 2378.170 ;
        RECT 571.630 2198.590 572.810 2199.770 ;
        RECT 573.230 2198.590 574.410 2199.770 ;
        RECT 571.630 2196.990 572.810 2198.170 ;
        RECT 573.230 2196.990 574.410 2198.170 ;
        RECT 571.630 2018.590 572.810 2019.770 ;
        RECT 573.230 2018.590 574.410 2019.770 ;
        RECT 571.630 2016.990 572.810 2018.170 ;
        RECT 573.230 2016.990 574.410 2018.170 ;
        RECT 571.630 1838.590 572.810 1839.770 ;
        RECT 573.230 1838.590 574.410 1839.770 ;
        RECT 571.630 1836.990 572.810 1838.170 ;
        RECT 573.230 1836.990 574.410 1838.170 ;
        RECT 571.630 1658.590 572.810 1659.770 ;
        RECT 573.230 1658.590 574.410 1659.770 ;
        RECT 571.630 1656.990 572.810 1658.170 ;
        RECT 573.230 1656.990 574.410 1658.170 ;
        RECT 571.630 1478.590 572.810 1479.770 ;
        RECT 573.230 1478.590 574.410 1479.770 ;
        RECT 571.630 1476.990 572.810 1478.170 ;
        RECT 573.230 1476.990 574.410 1478.170 ;
        RECT 571.630 1298.590 572.810 1299.770 ;
        RECT 573.230 1298.590 574.410 1299.770 ;
        RECT 571.630 1296.990 572.810 1298.170 ;
        RECT 573.230 1296.990 574.410 1298.170 ;
        RECT 571.630 1118.590 572.810 1119.770 ;
        RECT 573.230 1118.590 574.410 1119.770 ;
        RECT 571.630 1116.990 572.810 1118.170 ;
        RECT 573.230 1116.990 574.410 1118.170 ;
        RECT 571.630 938.590 572.810 939.770 ;
        RECT 573.230 938.590 574.410 939.770 ;
        RECT 571.630 936.990 572.810 938.170 ;
        RECT 573.230 936.990 574.410 938.170 ;
        RECT 751.630 3527.810 752.810 3528.990 ;
        RECT 753.230 3527.810 754.410 3528.990 ;
        RECT 751.630 3526.210 752.810 3527.390 ;
        RECT 753.230 3526.210 754.410 3527.390 ;
        RECT 751.630 3458.590 752.810 3459.770 ;
        RECT 753.230 3458.590 754.410 3459.770 ;
        RECT 751.630 3456.990 752.810 3458.170 ;
        RECT 753.230 3456.990 754.410 3458.170 ;
        RECT 751.630 3278.590 752.810 3279.770 ;
        RECT 753.230 3278.590 754.410 3279.770 ;
        RECT 751.630 3276.990 752.810 3278.170 ;
        RECT 753.230 3276.990 754.410 3278.170 ;
        RECT 751.630 3098.590 752.810 3099.770 ;
        RECT 753.230 3098.590 754.410 3099.770 ;
        RECT 751.630 3096.990 752.810 3098.170 ;
        RECT 753.230 3096.990 754.410 3098.170 ;
        RECT 751.630 2918.590 752.810 2919.770 ;
        RECT 753.230 2918.590 754.410 2919.770 ;
        RECT 751.630 2916.990 752.810 2918.170 ;
        RECT 753.230 2916.990 754.410 2918.170 ;
        RECT 751.630 2738.590 752.810 2739.770 ;
        RECT 753.230 2738.590 754.410 2739.770 ;
        RECT 751.630 2736.990 752.810 2738.170 ;
        RECT 753.230 2736.990 754.410 2738.170 ;
        RECT 751.630 2558.590 752.810 2559.770 ;
        RECT 753.230 2558.590 754.410 2559.770 ;
        RECT 751.630 2556.990 752.810 2558.170 ;
        RECT 753.230 2556.990 754.410 2558.170 ;
        RECT 751.630 2378.590 752.810 2379.770 ;
        RECT 753.230 2378.590 754.410 2379.770 ;
        RECT 751.630 2376.990 752.810 2378.170 ;
        RECT 753.230 2376.990 754.410 2378.170 ;
        RECT 751.630 2198.590 752.810 2199.770 ;
        RECT 753.230 2198.590 754.410 2199.770 ;
        RECT 751.630 2196.990 752.810 2198.170 ;
        RECT 753.230 2196.990 754.410 2198.170 ;
        RECT 751.630 2018.590 752.810 2019.770 ;
        RECT 753.230 2018.590 754.410 2019.770 ;
        RECT 751.630 2016.990 752.810 2018.170 ;
        RECT 753.230 2016.990 754.410 2018.170 ;
        RECT 751.630 1838.590 752.810 1839.770 ;
        RECT 753.230 1838.590 754.410 1839.770 ;
        RECT 751.630 1836.990 752.810 1838.170 ;
        RECT 753.230 1836.990 754.410 1838.170 ;
        RECT 751.630 1658.590 752.810 1659.770 ;
        RECT 753.230 1658.590 754.410 1659.770 ;
        RECT 751.630 1656.990 752.810 1658.170 ;
        RECT 753.230 1656.990 754.410 1658.170 ;
        RECT 751.630 1478.590 752.810 1479.770 ;
        RECT 753.230 1478.590 754.410 1479.770 ;
        RECT 751.630 1476.990 752.810 1478.170 ;
        RECT 753.230 1476.990 754.410 1478.170 ;
        RECT 751.630 1298.590 752.810 1299.770 ;
        RECT 753.230 1298.590 754.410 1299.770 ;
        RECT 751.630 1296.990 752.810 1298.170 ;
        RECT 753.230 1296.990 754.410 1298.170 ;
        RECT 751.630 1118.590 752.810 1119.770 ;
        RECT 753.230 1118.590 754.410 1119.770 ;
        RECT 751.630 1116.990 752.810 1118.170 ;
        RECT 753.230 1116.990 754.410 1118.170 ;
        RECT 751.630 938.590 752.810 939.770 ;
        RECT 753.230 938.590 754.410 939.770 ;
        RECT 751.630 936.990 752.810 938.170 ;
        RECT 753.230 936.990 754.410 938.170 ;
        RECT 211.630 758.590 212.810 759.770 ;
        RECT 213.230 758.590 214.410 759.770 ;
        RECT 211.630 756.990 212.810 758.170 ;
        RECT 213.230 756.990 214.410 758.170 ;
        RECT 211.630 578.590 212.810 579.770 ;
        RECT 213.230 578.590 214.410 579.770 ;
        RECT 211.630 576.990 212.810 578.170 ;
        RECT 213.230 576.990 214.410 578.170 ;
        RECT 498.050 758.590 499.230 759.770 ;
        RECT 498.050 756.990 499.230 758.170 ;
        RECT 498.050 578.590 499.230 579.770 ;
        RECT 498.050 576.990 499.230 578.170 ;
        RECT 651.650 758.590 652.830 759.770 ;
        RECT 651.650 756.990 652.830 758.170 ;
        RECT 651.650 578.590 652.830 579.770 ;
        RECT 651.650 576.990 652.830 578.170 ;
        RECT 751.630 758.590 752.810 759.770 ;
        RECT 753.230 758.590 754.410 759.770 ;
        RECT 751.630 756.990 752.810 758.170 ;
        RECT 753.230 756.990 754.410 758.170 ;
        RECT 751.630 578.590 752.810 579.770 ;
        RECT 753.230 578.590 754.410 579.770 ;
        RECT 751.630 576.990 752.810 578.170 ;
        RECT 753.230 576.990 754.410 578.170 ;
        RECT 211.630 398.590 212.810 399.770 ;
        RECT 213.230 398.590 214.410 399.770 ;
        RECT 211.630 396.990 212.810 398.170 ;
        RECT 213.230 396.990 214.410 398.170 ;
        RECT 211.630 218.590 212.810 219.770 ;
        RECT 213.230 218.590 214.410 219.770 ;
        RECT 211.630 216.990 212.810 218.170 ;
        RECT 213.230 216.990 214.410 218.170 ;
        RECT 211.630 38.590 212.810 39.770 ;
        RECT 213.230 38.590 214.410 39.770 ;
        RECT 211.630 36.990 212.810 38.170 ;
        RECT 213.230 36.990 214.410 38.170 ;
        RECT 211.630 -7.710 212.810 -6.530 ;
        RECT 213.230 -7.710 214.410 -6.530 ;
        RECT 211.630 -9.310 212.810 -8.130 ;
        RECT 213.230 -9.310 214.410 -8.130 ;
        RECT 391.630 398.590 392.810 399.770 ;
        RECT 393.230 398.590 394.410 399.770 ;
        RECT 391.630 396.990 392.810 398.170 ;
        RECT 393.230 396.990 394.410 398.170 ;
        RECT 391.630 218.590 392.810 219.770 ;
        RECT 393.230 218.590 394.410 219.770 ;
        RECT 391.630 216.990 392.810 218.170 ;
        RECT 393.230 216.990 394.410 218.170 ;
        RECT 391.630 38.590 392.810 39.770 ;
        RECT 393.230 38.590 394.410 39.770 ;
        RECT 391.630 36.990 392.810 38.170 ;
        RECT 393.230 36.990 394.410 38.170 ;
        RECT 391.630 -7.710 392.810 -6.530 ;
        RECT 393.230 -7.710 394.410 -6.530 ;
        RECT 391.630 -9.310 392.810 -8.130 ;
        RECT 393.230 -9.310 394.410 -8.130 ;
        RECT 571.630 398.590 572.810 399.770 ;
        RECT 573.230 398.590 574.410 399.770 ;
        RECT 571.630 396.990 572.810 398.170 ;
        RECT 573.230 396.990 574.410 398.170 ;
        RECT 571.630 218.590 572.810 219.770 ;
        RECT 573.230 218.590 574.410 219.770 ;
        RECT 571.630 216.990 572.810 218.170 ;
        RECT 573.230 216.990 574.410 218.170 ;
        RECT 571.630 38.590 572.810 39.770 ;
        RECT 573.230 38.590 574.410 39.770 ;
        RECT 571.630 36.990 572.810 38.170 ;
        RECT 573.230 36.990 574.410 38.170 ;
        RECT 571.630 -7.710 572.810 -6.530 ;
        RECT 573.230 -7.710 574.410 -6.530 ;
        RECT 571.630 -9.310 572.810 -8.130 ;
        RECT 573.230 -9.310 574.410 -8.130 ;
        RECT 751.630 398.590 752.810 399.770 ;
        RECT 753.230 398.590 754.410 399.770 ;
        RECT 751.630 396.990 752.810 398.170 ;
        RECT 753.230 396.990 754.410 398.170 ;
        RECT 751.630 218.590 752.810 219.770 ;
        RECT 753.230 218.590 754.410 219.770 ;
        RECT 751.630 216.990 752.810 218.170 ;
        RECT 753.230 216.990 754.410 218.170 ;
        RECT 751.630 38.590 752.810 39.770 ;
        RECT 753.230 38.590 754.410 39.770 ;
        RECT 751.630 36.990 752.810 38.170 ;
        RECT 753.230 36.990 754.410 38.170 ;
        RECT 751.630 -7.710 752.810 -6.530 ;
        RECT 753.230 -7.710 754.410 -6.530 ;
        RECT 751.630 -9.310 752.810 -8.130 ;
        RECT 753.230 -9.310 754.410 -8.130 ;
        RECT 931.630 3527.810 932.810 3528.990 ;
        RECT 933.230 3527.810 934.410 3528.990 ;
        RECT 931.630 3526.210 932.810 3527.390 ;
        RECT 933.230 3526.210 934.410 3527.390 ;
        RECT 931.630 3458.590 932.810 3459.770 ;
        RECT 933.230 3458.590 934.410 3459.770 ;
        RECT 931.630 3456.990 932.810 3458.170 ;
        RECT 933.230 3456.990 934.410 3458.170 ;
        RECT 931.630 3278.590 932.810 3279.770 ;
        RECT 933.230 3278.590 934.410 3279.770 ;
        RECT 931.630 3276.990 932.810 3278.170 ;
        RECT 933.230 3276.990 934.410 3278.170 ;
        RECT 931.630 3098.590 932.810 3099.770 ;
        RECT 933.230 3098.590 934.410 3099.770 ;
        RECT 931.630 3096.990 932.810 3098.170 ;
        RECT 933.230 3096.990 934.410 3098.170 ;
        RECT 931.630 2918.590 932.810 2919.770 ;
        RECT 933.230 2918.590 934.410 2919.770 ;
        RECT 931.630 2916.990 932.810 2918.170 ;
        RECT 933.230 2916.990 934.410 2918.170 ;
        RECT 931.630 2738.590 932.810 2739.770 ;
        RECT 933.230 2738.590 934.410 2739.770 ;
        RECT 931.630 2736.990 932.810 2738.170 ;
        RECT 933.230 2736.990 934.410 2738.170 ;
        RECT 931.630 2558.590 932.810 2559.770 ;
        RECT 933.230 2558.590 934.410 2559.770 ;
        RECT 931.630 2556.990 932.810 2558.170 ;
        RECT 933.230 2556.990 934.410 2558.170 ;
        RECT 931.630 2378.590 932.810 2379.770 ;
        RECT 933.230 2378.590 934.410 2379.770 ;
        RECT 931.630 2376.990 932.810 2378.170 ;
        RECT 933.230 2376.990 934.410 2378.170 ;
        RECT 931.630 2198.590 932.810 2199.770 ;
        RECT 933.230 2198.590 934.410 2199.770 ;
        RECT 931.630 2196.990 932.810 2198.170 ;
        RECT 933.230 2196.990 934.410 2198.170 ;
        RECT 931.630 2018.590 932.810 2019.770 ;
        RECT 933.230 2018.590 934.410 2019.770 ;
        RECT 931.630 2016.990 932.810 2018.170 ;
        RECT 933.230 2016.990 934.410 2018.170 ;
        RECT 931.630 1838.590 932.810 1839.770 ;
        RECT 933.230 1838.590 934.410 1839.770 ;
        RECT 931.630 1836.990 932.810 1838.170 ;
        RECT 933.230 1836.990 934.410 1838.170 ;
        RECT 931.630 1658.590 932.810 1659.770 ;
        RECT 933.230 1658.590 934.410 1659.770 ;
        RECT 931.630 1656.990 932.810 1658.170 ;
        RECT 933.230 1656.990 934.410 1658.170 ;
        RECT 931.630 1478.590 932.810 1479.770 ;
        RECT 933.230 1478.590 934.410 1479.770 ;
        RECT 931.630 1476.990 932.810 1478.170 ;
        RECT 933.230 1476.990 934.410 1478.170 ;
        RECT 931.630 1298.590 932.810 1299.770 ;
        RECT 933.230 1298.590 934.410 1299.770 ;
        RECT 931.630 1296.990 932.810 1298.170 ;
        RECT 933.230 1296.990 934.410 1298.170 ;
        RECT 931.630 1118.590 932.810 1119.770 ;
        RECT 933.230 1118.590 934.410 1119.770 ;
        RECT 931.630 1116.990 932.810 1118.170 ;
        RECT 933.230 1116.990 934.410 1118.170 ;
        RECT 931.630 938.590 932.810 939.770 ;
        RECT 933.230 938.590 934.410 939.770 ;
        RECT 931.630 936.990 932.810 938.170 ;
        RECT 933.230 936.990 934.410 938.170 ;
        RECT 931.630 758.590 932.810 759.770 ;
        RECT 933.230 758.590 934.410 759.770 ;
        RECT 931.630 756.990 932.810 758.170 ;
        RECT 933.230 756.990 934.410 758.170 ;
        RECT 931.630 578.590 932.810 579.770 ;
        RECT 933.230 578.590 934.410 579.770 ;
        RECT 931.630 576.990 932.810 578.170 ;
        RECT 933.230 576.990 934.410 578.170 ;
        RECT 931.630 398.590 932.810 399.770 ;
        RECT 933.230 398.590 934.410 399.770 ;
        RECT 931.630 396.990 932.810 398.170 ;
        RECT 933.230 396.990 934.410 398.170 ;
        RECT 931.630 218.590 932.810 219.770 ;
        RECT 933.230 218.590 934.410 219.770 ;
        RECT 931.630 216.990 932.810 218.170 ;
        RECT 933.230 216.990 934.410 218.170 ;
        RECT 931.630 38.590 932.810 39.770 ;
        RECT 933.230 38.590 934.410 39.770 ;
        RECT 931.630 36.990 932.810 38.170 ;
        RECT 933.230 36.990 934.410 38.170 ;
        RECT 931.630 -7.710 932.810 -6.530 ;
        RECT 933.230 -7.710 934.410 -6.530 ;
        RECT 931.630 -9.310 932.810 -8.130 ;
        RECT 933.230 -9.310 934.410 -8.130 ;
        RECT 1111.630 3527.810 1112.810 3528.990 ;
        RECT 1113.230 3527.810 1114.410 3528.990 ;
        RECT 1111.630 3526.210 1112.810 3527.390 ;
        RECT 1113.230 3526.210 1114.410 3527.390 ;
        RECT 1111.630 3458.590 1112.810 3459.770 ;
        RECT 1113.230 3458.590 1114.410 3459.770 ;
        RECT 1111.630 3456.990 1112.810 3458.170 ;
        RECT 1113.230 3456.990 1114.410 3458.170 ;
        RECT 1111.630 3278.590 1112.810 3279.770 ;
        RECT 1113.230 3278.590 1114.410 3279.770 ;
        RECT 1111.630 3276.990 1112.810 3278.170 ;
        RECT 1113.230 3276.990 1114.410 3278.170 ;
        RECT 1111.630 3098.590 1112.810 3099.770 ;
        RECT 1113.230 3098.590 1114.410 3099.770 ;
        RECT 1111.630 3096.990 1112.810 3098.170 ;
        RECT 1113.230 3096.990 1114.410 3098.170 ;
        RECT 1111.630 2918.590 1112.810 2919.770 ;
        RECT 1113.230 2918.590 1114.410 2919.770 ;
        RECT 1111.630 2916.990 1112.810 2918.170 ;
        RECT 1113.230 2916.990 1114.410 2918.170 ;
        RECT 1111.630 2738.590 1112.810 2739.770 ;
        RECT 1113.230 2738.590 1114.410 2739.770 ;
        RECT 1111.630 2736.990 1112.810 2738.170 ;
        RECT 1113.230 2736.990 1114.410 2738.170 ;
        RECT 1111.630 2558.590 1112.810 2559.770 ;
        RECT 1113.230 2558.590 1114.410 2559.770 ;
        RECT 1111.630 2556.990 1112.810 2558.170 ;
        RECT 1113.230 2556.990 1114.410 2558.170 ;
        RECT 1111.630 2378.590 1112.810 2379.770 ;
        RECT 1113.230 2378.590 1114.410 2379.770 ;
        RECT 1111.630 2376.990 1112.810 2378.170 ;
        RECT 1113.230 2376.990 1114.410 2378.170 ;
        RECT 1111.630 2198.590 1112.810 2199.770 ;
        RECT 1113.230 2198.590 1114.410 2199.770 ;
        RECT 1111.630 2196.990 1112.810 2198.170 ;
        RECT 1113.230 2196.990 1114.410 2198.170 ;
        RECT 1111.630 2018.590 1112.810 2019.770 ;
        RECT 1113.230 2018.590 1114.410 2019.770 ;
        RECT 1111.630 2016.990 1112.810 2018.170 ;
        RECT 1113.230 2016.990 1114.410 2018.170 ;
        RECT 1111.630 1838.590 1112.810 1839.770 ;
        RECT 1113.230 1838.590 1114.410 1839.770 ;
        RECT 1111.630 1836.990 1112.810 1838.170 ;
        RECT 1113.230 1836.990 1114.410 1838.170 ;
        RECT 1111.630 1658.590 1112.810 1659.770 ;
        RECT 1113.230 1658.590 1114.410 1659.770 ;
        RECT 1111.630 1656.990 1112.810 1658.170 ;
        RECT 1113.230 1656.990 1114.410 1658.170 ;
        RECT 1111.630 1478.590 1112.810 1479.770 ;
        RECT 1113.230 1478.590 1114.410 1479.770 ;
        RECT 1111.630 1476.990 1112.810 1478.170 ;
        RECT 1113.230 1476.990 1114.410 1478.170 ;
        RECT 1111.630 1298.590 1112.810 1299.770 ;
        RECT 1113.230 1298.590 1114.410 1299.770 ;
        RECT 1111.630 1296.990 1112.810 1298.170 ;
        RECT 1113.230 1296.990 1114.410 1298.170 ;
        RECT 1111.630 1118.590 1112.810 1119.770 ;
        RECT 1113.230 1118.590 1114.410 1119.770 ;
        RECT 1111.630 1116.990 1112.810 1118.170 ;
        RECT 1113.230 1116.990 1114.410 1118.170 ;
        RECT 1111.630 938.590 1112.810 939.770 ;
        RECT 1113.230 938.590 1114.410 939.770 ;
        RECT 1111.630 936.990 1112.810 938.170 ;
        RECT 1113.230 936.990 1114.410 938.170 ;
        RECT 1111.630 758.590 1112.810 759.770 ;
        RECT 1113.230 758.590 1114.410 759.770 ;
        RECT 1111.630 756.990 1112.810 758.170 ;
        RECT 1113.230 756.990 1114.410 758.170 ;
        RECT 1111.630 578.590 1112.810 579.770 ;
        RECT 1113.230 578.590 1114.410 579.770 ;
        RECT 1111.630 576.990 1112.810 578.170 ;
        RECT 1113.230 576.990 1114.410 578.170 ;
        RECT 1111.630 398.590 1112.810 399.770 ;
        RECT 1113.230 398.590 1114.410 399.770 ;
        RECT 1111.630 396.990 1112.810 398.170 ;
        RECT 1113.230 396.990 1114.410 398.170 ;
        RECT 1111.630 218.590 1112.810 219.770 ;
        RECT 1113.230 218.590 1114.410 219.770 ;
        RECT 1111.630 216.990 1112.810 218.170 ;
        RECT 1113.230 216.990 1114.410 218.170 ;
        RECT 1111.630 38.590 1112.810 39.770 ;
        RECT 1113.230 38.590 1114.410 39.770 ;
        RECT 1111.630 36.990 1112.810 38.170 ;
        RECT 1113.230 36.990 1114.410 38.170 ;
        RECT 1111.630 -7.710 1112.810 -6.530 ;
        RECT 1113.230 -7.710 1114.410 -6.530 ;
        RECT 1111.630 -9.310 1112.810 -8.130 ;
        RECT 1113.230 -9.310 1114.410 -8.130 ;
        RECT 1291.630 3527.810 1292.810 3528.990 ;
        RECT 1293.230 3527.810 1294.410 3528.990 ;
        RECT 1291.630 3526.210 1292.810 3527.390 ;
        RECT 1293.230 3526.210 1294.410 3527.390 ;
        RECT 1291.630 3458.590 1292.810 3459.770 ;
        RECT 1293.230 3458.590 1294.410 3459.770 ;
        RECT 1291.630 3456.990 1292.810 3458.170 ;
        RECT 1293.230 3456.990 1294.410 3458.170 ;
        RECT 1291.630 3278.590 1292.810 3279.770 ;
        RECT 1293.230 3278.590 1294.410 3279.770 ;
        RECT 1291.630 3276.990 1292.810 3278.170 ;
        RECT 1293.230 3276.990 1294.410 3278.170 ;
        RECT 1291.630 3098.590 1292.810 3099.770 ;
        RECT 1293.230 3098.590 1294.410 3099.770 ;
        RECT 1291.630 3096.990 1292.810 3098.170 ;
        RECT 1293.230 3096.990 1294.410 3098.170 ;
        RECT 1291.630 2918.590 1292.810 2919.770 ;
        RECT 1293.230 2918.590 1294.410 2919.770 ;
        RECT 1291.630 2916.990 1292.810 2918.170 ;
        RECT 1293.230 2916.990 1294.410 2918.170 ;
        RECT 1291.630 2738.590 1292.810 2739.770 ;
        RECT 1293.230 2738.590 1294.410 2739.770 ;
        RECT 1291.630 2736.990 1292.810 2738.170 ;
        RECT 1293.230 2736.990 1294.410 2738.170 ;
        RECT 1291.630 2558.590 1292.810 2559.770 ;
        RECT 1293.230 2558.590 1294.410 2559.770 ;
        RECT 1291.630 2556.990 1292.810 2558.170 ;
        RECT 1293.230 2556.990 1294.410 2558.170 ;
        RECT 1291.630 2378.590 1292.810 2379.770 ;
        RECT 1293.230 2378.590 1294.410 2379.770 ;
        RECT 1291.630 2376.990 1292.810 2378.170 ;
        RECT 1293.230 2376.990 1294.410 2378.170 ;
        RECT 1291.630 2198.590 1292.810 2199.770 ;
        RECT 1293.230 2198.590 1294.410 2199.770 ;
        RECT 1291.630 2196.990 1292.810 2198.170 ;
        RECT 1293.230 2196.990 1294.410 2198.170 ;
        RECT 1291.630 2018.590 1292.810 2019.770 ;
        RECT 1293.230 2018.590 1294.410 2019.770 ;
        RECT 1291.630 2016.990 1292.810 2018.170 ;
        RECT 1293.230 2016.990 1294.410 2018.170 ;
        RECT 1291.630 1838.590 1292.810 1839.770 ;
        RECT 1293.230 1838.590 1294.410 1839.770 ;
        RECT 1291.630 1836.990 1292.810 1838.170 ;
        RECT 1293.230 1836.990 1294.410 1838.170 ;
        RECT 1291.630 1658.590 1292.810 1659.770 ;
        RECT 1293.230 1658.590 1294.410 1659.770 ;
        RECT 1291.630 1656.990 1292.810 1658.170 ;
        RECT 1293.230 1656.990 1294.410 1658.170 ;
        RECT 1291.630 1478.590 1292.810 1479.770 ;
        RECT 1293.230 1478.590 1294.410 1479.770 ;
        RECT 1291.630 1476.990 1292.810 1478.170 ;
        RECT 1293.230 1476.990 1294.410 1478.170 ;
        RECT 1291.630 1298.590 1292.810 1299.770 ;
        RECT 1293.230 1298.590 1294.410 1299.770 ;
        RECT 1291.630 1296.990 1292.810 1298.170 ;
        RECT 1293.230 1296.990 1294.410 1298.170 ;
        RECT 1291.630 1118.590 1292.810 1119.770 ;
        RECT 1293.230 1118.590 1294.410 1119.770 ;
        RECT 1291.630 1116.990 1292.810 1118.170 ;
        RECT 1293.230 1116.990 1294.410 1118.170 ;
        RECT 1291.630 938.590 1292.810 939.770 ;
        RECT 1293.230 938.590 1294.410 939.770 ;
        RECT 1291.630 936.990 1292.810 938.170 ;
        RECT 1293.230 936.990 1294.410 938.170 ;
        RECT 1291.630 758.590 1292.810 759.770 ;
        RECT 1293.230 758.590 1294.410 759.770 ;
        RECT 1291.630 756.990 1292.810 758.170 ;
        RECT 1293.230 756.990 1294.410 758.170 ;
        RECT 1291.630 578.590 1292.810 579.770 ;
        RECT 1293.230 578.590 1294.410 579.770 ;
        RECT 1291.630 576.990 1292.810 578.170 ;
        RECT 1293.230 576.990 1294.410 578.170 ;
        RECT 1291.630 398.590 1292.810 399.770 ;
        RECT 1293.230 398.590 1294.410 399.770 ;
        RECT 1291.630 396.990 1292.810 398.170 ;
        RECT 1293.230 396.990 1294.410 398.170 ;
        RECT 1291.630 218.590 1292.810 219.770 ;
        RECT 1293.230 218.590 1294.410 219.770 ;
        RECT 1291.630 216.990 1292.810 218.170 ;
        RECT 1293.230 216.990 1294.410 218.170 ;
        RECT 1291.630 38.590 1292.810 39.770 ;
        RECT 1293.230 38.590 1294.410 39.770 ;
        RECT 1291.630 36.990 1292.810 38.170 ;
        RECT 1293.230 36.990 1294.410 38.170 ;
        RECT 1291.630 -7.710 1292.810 -6.530 ;
        RECT 1293.230 -7.710 1294.410 -6.530 ;
        RECT 1291.630 -9.310 1292.810 -8.130 ;
        RECT 1293.230 -9.310 1294.410 -8.130 ;
        RECT 1471.630 3527.810 1472.810 3528.990 ;
        RECT 1473.230 3527.810 1474.410 3528.990 ;
        RECT 1471.630 3526.210 1472.810 3527.390 ;
        RECT 1473.230 3526.210 1474.410 3527.390 ;
        RECT 1471.630 3458.590 1472.810 3459.770 ;
        RECT 1473.230 3458.590 1474.410 3459.770 ;
        RECT 1471.630 3456.990 1472.810 3458.170 ;
        RECT 1473.230 3456.990 1474.410 3458.170 ;
        RECT 1471.630 3278.590 1472.810 3279.770 ;
        RECT 1473.230 3278.590 1474.410 3279.770 ;
        RECT 1471.630 3276.990 1472.810 3278.170 ;
        RECT 1473.230 3276.990 1474.410 3278.170 ;
        RECT 1471.630 3098.590 1472.810 3099.770 ;
        RECT 1473.230 3098.590 1474.410 3099.770 ;
        RECT 1471.630 3096.990 1472.810 3098.170 ;
        RECT 1473.230 3096.990 1474.410 3098.170 ;
        RECT 1471.630 2918.590 1472.810 2919.770 ;
        RECT 1473.230 2918.590 1474.410 2919.770 ;
        RECT 1471.630 2916.990 1472.810 2918.170 ;
        RECT 1473.230 2916.990 1474.410 2918.170 ;
        RECT 1471.630 2738.590 1472.810 2739.770 ;
        RECT 1473.230 2738.590 1474.410 2739.770 ;
        RECT 1471.630 2736.990 1472.810 2738.170 ;
        RECT 1473.230 2736.990 1474.410 2738.170 ;
        RECT 1471.630 2558.590 1472.810 2559.770 ;
        RECT 1473.230 2558.590 1474.410 2559.770 ;
        RECT 1471.630 2556.990 1472.810 2558.170 ;
        RECT 1473.230 2556.990 1474.410 2558.170 ;
        RECT 1471.630 2378.590 1472.810 2379.770 ;
        RECT 1473.230 2378.590 1474.410 2379.770 ;
        RECT 1471.630 2376.990 1472.810 2378.170 ;
        RECT 1473.230 2376.990 1474.410 2378.170 ;
        RECT 1471.630 2198.590 1472.810 2199.770 ;
        RECT 1473.230 2198.590 1474.410 2199.770 ;
        RECT 1471.630 2196.990 1472.810 2198.170 ;
        RECT 1473.230 2196.990 1474.410 2198.170 ;
        RECT 1471.630 2018.590 1472.810 2019.770 ;
        RECT 1473.230 2018.590 1474.410 2019.770 ;
        RECT 1471.630 2016.990 1472.810 2018.170 ;
        RECT 1473.230 2016.990 1474.410 2018.170 ;
        RECT 1471.630 1838.590 1472.810 1839.770 ;
        RECT 1473.230 1838.590 1474.410 1839.770 ;
        RECT 1471.630 1836.990 1472.810 1838.170 ;
        RECT 1473.230 1836.990 1474.410 1838.170 ;
        RECT 1471.630 1658.590 1472.810 1659.770 ;
        RECT 1473.230 1658.590 1474.410 1659.770 ;
        RECT 1471.630 1656.990 1472.810 1658.170 ;
        RECT 1473.230 1656.990 1474.410 1658.170 ;
        RECT 1471.630 1478.590 1472.810 1479.770 ;
        RECT 1473.230 1478.590 1474.410 1479.770 ;
        RECT 1471.630 1476.990 1472.810 1478.170 ;
        RECT 1473.230 1476.990 1474.410 1478.170 ;
        RECT 1471.630 1298.590 1472.810 1299.770 ;
        RECT 1473.230 1298.590 1474.410 1299.770 ;
        RECT 1471.630 1296.990 1472.810 1298.170 ;
        RECT 1473.230 1296.990 1474.410 1298.170 ;
        RECT 1471.630 1118.590 1472.810 1119.770 ;
        RECT 1473.230 1118.590 1474.410 1119.770 ;
        RECT 1471.630 1116.990 1472.810 1118.170 ;
        RECT 1473.230 1116.990 1474.410 1118.170 ;
        RECT 1471.630 938.590 1472.810 939.770 ;
        RECT 1473.230 938.590 1474.410 939.770 ;
        RECT 1471.630 936.990 1472.810 938.170 ;
        RECT 1473.230 936.990 1474.410 938.170 ;
        RECT 1471.630 758.590 1472.810 759.770 ;
        RECT 1473.230 758.590 1474.410 759.770 ;
        RECT 1471.630 756.990 1472.810 758.170 ;
        RECT 1473.230 756.990 1474.410 758.170 ;
        RECT 1471.630 578.590 1472.810 579.770 ;
        RECT 1473.230 578.590 1474.410 579.770 ;
        RECT 1471.630 576.990 1472.810 578.170 ;
        RECT 1473.230 576.990 1474.410 578.170 ;
        RECT 1471.630 398.590 1472.810 399.770 ;
        RECT 1473.230 398.590 1474.410 399.770 ;
        RECT 1471.630 396.990 1472.810 398.170 ;
        RECT 1473.230 396.990 1474.410 398.170 ;
        RECT 1471.630 218.590 1472.810 219.770 ;
        RECT 1473.230 218.590 1474.410 219.770 ;
        RECT 1471.630 216.990 1472.810 218.170 ;
        RECT 1473.230 216.990 1474.410 218.170 ;
        RECT 1471.630 38.590 1472.810 39.770 ;
        RECT 1473.230 38.590 1474.410 39.770 ;
        RECT 1471.630 36.990 1472.810 38.170 ;
        RECT 1473.230 36.990 1474.410 38.170 ;
        RECT 1471.630 -7.710 1472.810 -6.530 ;
        RECT 1473.230 -7.710 1474.410 -6.530 ;
        RECT 1471.630 -9.310 1472.810 -8.130 ;
        RECT 1473.230 -9.310 1474.410 -8.130 ;
        RECT 1651.630 3527.810 1652.810 3528.990 ;
        RECT 1653.230 3527.810 1654.410 3528.990 ;
        RECT 1651.630 3526.210 1652.810 3527.390 ;
        RECT 1653.230 3526.210 1654.410 3527.390 ;
        RECT 1651.630 3458.590 1652.810 3459.770 ;
        RECT 1653.230 3458.590 1654.410 3459.770 ;
        RECT 1651.630 3456.990 1652.810 3458.170 ;
        RECT 1653.230 3456.990 1654.410 3458.170 ;
        RECT 1651.630 3278.590 1652.810 3279.770 ;
        RECT 1653.230 3278.590 1654.410 3279.770 ;
        RECT 1651.630 3276.990 1652.810 3278.170 ;
        RECT 1653.230 3276.990 1654.410 3278.170 ;
        RECT 1651.630 3098.590 1652.810 3099.770 ;
        RECT 1653.230 3098.590 1654.410 3099.770 ;
        RECT 1651.630 3096.990 1652.810 3098.170 ;
        RECT 1653.230 3096.990 1654.410 3098.170 ;
        RECT 1651.630 2918.590 1652.810 2919.770 ;
        RECT 1653.230 2918.590 1654.410 2919.770 ;
        RECT 1651.630 2916.990 1652.810 2918.170 ;
        RECT 1653.230 2916.990 1654.410 2918.170 ;
        RECT 1651.630 2738.590 1652.810 2739.770 ;
        RECT 1653.230 2738.590 1654.410 2739.770 ;
        RECT 1651.630 2736.990 1652.810 2738.170 ;
        RECT 1653.230 2736.990 1654.410 2738.170 ;
        RECT 1651.630 2558.590 1652.810 2559.770 ;
        RECT 1653.230 2558.590 1654.410 2559.770 ;
        RECT 1651.630 2556.990 1652.810 2558.170 ;
        RECT 1653.230 2556.990 1654.410 2558.170 ;
        RECT 1651.630 2378.590 1652.810 2379.770 ;
        RECT 1653.230 2378.590 1654.410 2379.770 ;
        RECT 1651.630 2376.990 1652.810 2378.170 ;
        RECT 1653.230 2376.990 1654.410 2378.170 ;
        RECT 1651.630 2198.590 1652.810 2199.770 ;
        RECT 1653.230 2198.590 1654.410 2199.770 ;
        RECT 1651.630 2196.990 1652.810 2198.170 ;
        RECT 1653.230 2196.990 1654.410 2198.170 ;
        RECT 1651.630 2018.590 1652.810 2019.770 ;
        RECT 1653.230 2018.590 1654.410 2019.770 ;
        RECT 1651.630 2016.990 1652.810 2018.170 ;
        RECT 1653.230 2016.990 1654.410 2018.170 ;
        RECT 1651.630 1838.590 1652.810 1839.770 ;
        RECT 1653.230 1838.590 1654.410 1839.770 ;
        RECT 1651.630 1836.990 1652.810 1838.170 ;
        RECT 1653.230 1836.990 1654.410 1838.170 ;
        RECT 1651.630 1658.590 1652.810 1659.770 ;
        RECT 1653.230 1658.590 1654.410 1659.770 ;
        RECT 1651.630 1656.990 1652.810 1658.170 ;
        RECT 1653.230 1656.990 1654.410 1658.170 ;
        RECT 1651.630 1478.590 1652.810 1479.770 ;
        RECT 1653.230 1478.590 1654.410 1479.770 ;
        RECT 1651.630 1476.990 1652.810 1478.170 ;
        RECT 1653.230 1476.990 1654.410 1478.170 ;
        RECT 1651.630 1298.590 1652.810 1299.770 ;
        RECT 1653.230 1298.590 1654.410 1299.770 ;
        RECT 1651.630 1296.990 1652.810 1298.170 ;
        RECT 1653.230 1296.990 1654.410 1298.170 ;
        RECT 1651.630 1118.590 1652.810 1119.770 ;
        RECT 1653.230 1118.590 1654.410 1119.770 ;
        RECT 1651.630 1116.990 1652.810 1118.170 ;
        RECT 1653.230 1116.990 1654.410 1118.170 ;
        RECT 1651.630 938.590 1652.810 939.770 ;
        RECT 1653.230 938.590 1654.410 939.770 ;
        RECT 1651.630 936.990 1652.810 938.170 ;
        RECT 1653.230 936.990 1654.410 938.170 ;
        RECT 1651.630 758.590 1652.810 759.770 ;
        RECT 1653.230 758.590 1654.410 759.770 ;
        RECT 1651.630 756.990 1652.810 758.170 ;
        RECT 1653.230 756.990 1654.410 758.170 ;
        RECT 1651.630 578.590 1652.810 579.770 ;
        RECT 1653.230 578.590 1654.410 579.770 ;
        RECT 1651.630 576.990 1652.810 578.170 ;
        RECT 1653.230 576.990 1654.410 578.170 ;
        RECT 1651.630 398.590 1652.810 399.770 ;
        RECT 1653.230 398.590 1654.410 399.770 ;
        RECT 1651.630 396.990 1652.810 398.170 ;
        RECT 1653.230 396.990 1654.410 398.170 ;
        RECT 1651.630 218.590 1652.810 219.770 ;
        RECT 1653.230 218.590 1654.410 219.770 ;
        RECT 1651.630 216.990 1652.810 218.170 ;
        RECT 1653.230 216.990 1654.410 218.170 ;
        RECT 1651.630 38.590 1652.810 39.770 ;
        RECT 1653.230 38.590 1654.410 39.770 ;
        RECT 1651.630 36.990 1652.810 38.170 ;
        RECT 1653.230 36.990 1654.410 38.170 ;
        RECT 1651.630 -7.710 1652.810 -6.530 ;
        RECT 1653.230 -7.710 1654.410 -6.530 ;
        RECT 1651.630 -9.310 1652.810 -8.130 ;
        RECT 1653.230 -9.310 1654.410 -8.130 ;
        RECT 1831.630 3527.810 1832.810 3528.990 ;
        RECT 1833.230 3527.810 1834.410 3528.990 ;
        RECT 1831.630 3526.210 1832.810 3527.390 ;
        RECT 1833.230 3526.210 1834.410 3527.390 ;
        RECT 1831.630 3458.590 1832.810 3459.770 ;
        RECT 1833.230 3458.590 1834.410 3459.770 ;
        RECT 1831.630 3456.990 1832.810 3458.170 ;
        RECT 1833.230 3456.990 1834.410 3458.170 ;
        RECT 1831.630 3278.590 1832.810 3279.770 ;
        RECT 1833.230 3278.590 1834.410 3279.770 ;
        RECT 1831.630 3276.990 1832.810 3278.170 ;
        RECT 1833.230 3276.990 1834.410 3278.170 ;
        RECT 1831.630 3098.590 1832.810 3099.770 ;
        RECT 1833.230 3098.590 1834.410 3099.770 ;
        RECT 1831.630 3096.990 1832.810 3098.170 ;
        RECT 1833.230 3096.990 1834.410 3098.170 ;
        RECT 1831.630 2918.590 1832.810 2919.770 ;
        RECT 1833.230 2918.590 1834.410 2919.770 ;
        RECT 1831.630 2916.990 1832.810 2918.170 ;
        RECT 1833.230 2916.990 1834.410 2918.170 ;
        RECT 1831.630 2738.590 1832.810 2739.770 ;
        RECT 1833.230 2738.590 1834.410 2739.770 ;
        RECT 1831.630 2736.990 1832.810 2738.170 ;
        RECT 1833.230 2736.990 1834.410 2738.170 ;
        RECT 1831.630 2558.590 1832.810 2559.770 ;
        RECT 1833.230 2558.590 1834.410 2559.770 ;
        RECT 1831.630 2556.990 1832.810 2558.170 ;
        RECT 1833.230 2556.990 1834.410 2558.170 ;
        RECT 1831.630 2378.590 1832.810 2379.770 ;
        RECT 1833.230 2378.590 1834.410 2379.770 ;
        RECT 1831.630 2376.990 1832.810 2378.170 ;
        RECT 1833.230 2376.990 1834.410 2378.170 ;
        RECT 1831.630 2198.590 1832.810 2199.770 ;
        RECT 1833.230 2198.590 1834.410 2199.770 ;
        RECT 1831.630 2196.990 1832.810 2198.170 ;
        RECT 1833.230 2196.990 1834.410 2198.170 ;
        RECT 1831.630 2018.590 1832.810 2019.770 ;
        RECT 1833.230 2018.590 1834.410 2019.770 ;
        RECT 1831.630 2016.990 1832.810 2018.170 ;
        RECT 1833.230 2016.990 1834.410 2018.170 ;
        RECT 1831.630 1838.590 1832.810 1839.770 ;
        RECT 1833.230 1838.590 1834.410 1839.770 ;
        RECT 1831.630 1836.990 1832.810 1838.170 ;
        RECT 1833.230 1836.990 1834.410 1838.170 ;
        RECT 1831.630 1658.590 1832.810 1659.770 ;
        RECT 1833.230 1658.590 1834.410 1659.770 ;
        RECT 1831.630 1656.990 1832.810 1658.170 ;
        RECT 1833.230 1656.990 1834.410 1658.170 ;
        RECT 1831.630 1478.590 1832.810 1479.770 ;
        RECT 1833.230 1478.590 1834.410 1479.770 ;
        RECT 1831.630 1476.990 1832.810 1478.170 ;
        RECT 1833.230 1476.990 1834.410 1478.170 ;
        RECT 1831.630 1298.590 1832.810 1299.770 ;
        RECT 1833.230 1298.590 1834.410 1299.770 ;
        RECT 1831.630 1296.990 1832.810 1298.170 ;
        RECT 1833.230 1296.990 1834.410 1298.170 ;
        RECT 1831.630 1118.590 1832.810 1119.770 ;
        RECT 1833.230 1118.590 1834.410 1119.770 ;
        RECT 1831.630 1116.990 1832.810 1118.170 ;
        RECT 1833.230 1116.990 1834.410 1118.170 ;
        RECT 1831.630 938.590 1832.810 939.770 ;
        RECT 1833.230 938.590 1834.410 939.770 ;
        RECT 1831.630 936.990 1832.810 938.170 ;
        RECT 1833.230 936.990 1834.410 938.170 ;
        RECT 1831.630 758.590 1832.810 759.770 ;
        RECT 1833.230 758.590 1834.410 759.770 ;
        RECT 1831.630 756.990 1832.810 758.170 ;
        RECT 1833.230 756.990 1834.410 758.170 ;
        RECT 1831.630 578.590 1832.810 579.770 ;
        RECT 1833.230 578.590 1834.410 579.770 ;
        RECT 1831.630 576.990 1832.810 578.170 ;
        RECT 1833.230 576.990 1834.410 578.170 ;
        RECT 1831.630 398.590 1832.810 399.770 ;
        RECT 1833.230 398.590 1834.410 399.770 ;
        RECT 1831.630 396.990 1832.810 398.170 ;
        RECT 1833.230 396.990 1834.410 398.170 ;
        RECT 1831.630 218.590 1832.810 219.770 ;
        RECT 1833.230 218.590 1834.410 219.770 ;
        RECT 1831.630 216.990 1832.810 218.170 ;
        RECT 1833.230 216.990 1834.410 218.170 ;
        RECT 1831.630 38.590 1832.810 39.770 ;
        RECT 1833.230 38.590 1834.410 39.770 ;
        RECT 1831.630 36.990 1832.810 38.170 ;
        RECT 1833.230 36.990 1834.410 38.170 ;
        RECT 1831.630 -7.710 1832.810 -6.530 ;
        RECT 1833.230 -7.710 1834.410 -6.530 ;
        RECT 1831.630 -9.310 1832.810 -8.130 ;
        RECT 1833.230 -9.310 1834.410 -8.130 ;
        RECT 2011.630 3527.810 2012.810 3528.990 ;
        RECT 2013.230 3527.810 2014.410 3528.990 ;
        RECT 2011.630 3526.210 2012.810 3527.390 ;
        RECT 2013.230 3526.210 2014.410 3527.390 ;
        RECT 2011.630 3458.590 2012.810 3459.770 ;
        RECT 2013.230 3458.590 2014.410 3459.770 ;
        RECT 2011.630 3456.990 2012.810 3458.170 ;
        RECT 2013.230 3456.990 2014.410 3458.170 ;
        RECT 2011.630 3278.590 2012.810 3279.770 ;
        RECT 2013.230 3278.590 2014.410 3279.770 ;
        RECT 2011.630 3276.990 2012.810 3278.170 ;
        RECT 2013.230 3276.990 2014.410 3278.170 ;
        RECT 2011.630 3098.590 2012.810 3099.770 ;
        RECT 2013.230 3098.590 2014.410 3099.770 ;
        RECT 2011.630 3096.990 2012.810 3098.170 ;
        RECT 2013.230 3096.990 2014.410 3098.170 ;
        RECT 2011.630 2918.590 2012.810 2919.770 ;
        RECT 2013.230 2918.590 2014.410 2919.770 ;
        RECT 2011.630 2916.990 2012.810 2918.170 ;
        RECT 2013.230 2916.990 2014.410 2918.170 ;
        RECT 2011.630 2738.590 2012.810 2739.770 ;
        RECT 2013.230 2738.590 2014.410 2739.770 ;
        RECT 2011.630 2736.990 2012.810 2738.170 ;
        RECT 2013.230 2736.990 2014.410 2738.170 ;
        RECT 2011.630 2558.590 2012.810 2559.770 ;
        RECT 2013.230 2558.590 2014.410 2559.770 ;
        RECT 2011.630 2556.990 2012.810 2558.170 ;
        RECT 2013.230 2556.990 2014.410 2558.170 ;
        RECT 2011.630 2378.590 2012.810 2379.770 ;
        RECT 2013.230 2378.590 2014.410 2379.770 ;
        RECT 2011.630 2376.990 2012.810 2378.170 ;
        RECT 2013.230 2376.990 2014.410 2378.170 ;
        RECT 2011.630 2198.590 2012.810 2199.770 ;
        RECT 2013.230 2198.590 2014.410 2199.770 ;
        RECT 2011.630 2196.990 2012.810 2198.170 ;
        RECT 2013.230 2196.990 2014.410 2198.170 ;
        RECT 2011.630 2018.590 2012.810 2019.770 ;
        RECT 2013.230 2018.590 2014.410 2019.770 ;
        RECT 2011.630 2016.990 2012.810 2018.170 ;
        RECT 2013.230 2016.990 2014.410 2018.170 ;
        RECT 2011.630 1838.590 2012.810 1839.770 ;
        RECT 2013.230 1838.590 2014.410 1839.770 ;
        RECT 2011.630 1836.990 2012.810 1838.170 ;
        RECT 2013.230 1836.990 2014.410 1838.170 ;
        RECT 2011.630 1658.590 2012.810 1659.770 ;
        RECT 2013.230 1658.590 2014.410 1659.770 ;
        RECT 2011.630 1656.990 2012.810 1658.170 ;
        RECT 2013.230 1656.990 2014.410 1658.170 ;
        RECT 2011.630 1478.590 2012.810 1479.770 ;
        RECT 2013.230 1478.590 2014.410 1479.770 ;
        RECT 2011.630 1476.990 2012.810 1478.170 ;
        RECT 2013.230 1476.990 2014.410 1478.170 ;
        RECT 2011.630 1298.590 2012.810 1299.770 ;
        RECT 2013.230 1298.590 2014.410 1299.770 ;
        RECT 2011.630 1296.990 2012.810 1298.170 ;
        RECT 2013.230 1296.990 2014.410 1298.170 ;
        RECT 2011.630 1118.590 2012.810 1119.770 ;
        RECT 2013.230 1118.590 2014.410 1119.770 ;
        RECT 2011.630 1116.990 2012.810 1118.170 ;
        RECT 2013.230 1116.990 2014.410 1118.170 ;
        RECT 2011.630 938.590 2012.810 939.770 ;
        RECT 2013.230 938.590 2014.410 939.770 ;
        RECT 2011.630 936.990 2012.810 938.170 ;
        RECT 2013.230 936.990 2014.410 938.170 ;
        RECT 2011.630 758.590 2012.810 759.770 ;
        RECT 2013.230 758.590 2014.410 759.770 ;
        RECT 2011.630 756.990 2012.810 758.170 ;
        RECT 2013.230 756.990 2014.410 758.170 ;
        RECT 2011.630 578.590 2012.810 579.770 ;
        RECT 2013.230 578.590 2014.410 579.770 ;
        RECT 2011.630 576.990 2012.810 578.170 ;
        RECT 2013.230 576.990 2014.410 578.170 ;
        RECT 2011.630 398.590 2012.810 399.770 ;
        RECT 2013.230 398.590 2014.410 399.770 ;
        RECT 2011.630 396.990 2012.810 398.170 ;
        RECT 2013.230 396.990 2014.410 398.170 ;
        RECT 2011.630 218.590 2012.810 219.770 ;
        RECT 2013.230 218.590 2014.410 219.770 ;
        RECT 2011.630 216.990 2012.810 218.170 ;
        RECT 2013.230 216.990 2014.410 218.170 ;
        RECT 2011.630 38.590 2012.810 39.770 ;
        RECT 2013.230 38.590 2014.410 39.770 ;
        RECT 2011.630 36.990 2012.810 38.170 ;
        RECT 2013.230 36.990 2014.410 38.170 ;
        RECT 2011.630 -7.710 2012.810 -6.530 ;
        RECT 2013.230 -7.710 2014.410 -6.530 ;
        RECT 2011.630 -9.310 2012.810 -8.130 ;
        RECT 2013.230 -9.310 2014.410 -8.130 ;
        RECT 2191.630 3527.810 2192.810 3528.990 ;
        RECT 2193.230 3527.810 2194.410 3528.990 ;
        RECT 2191.630 3526.210 2192.810 3527.390 ;
        RECT 2193.230 3526.210 2194.410 3527.390 ;
        RECT 2191.630 3458.590 2192.810 3459.770 ;
        RECT 2193.230 3458.590 2194.410 3459.770 ;
        RECT 2191.630 3456.990 2192.810 3458.170 ;
        RECT 2193.230 3456.990 2194.410 3458.170 ;
        RECT 2191.630 3278.590 2192.810 3279.770 ;
        RECT 2193.230 3278.590 2194.410 3279.770 ;
        RECT 2191.630 3276.990 2192.810 3278.170 ;
        RECT 2193.230 3276.990 2194.410 3278.170 ;
        RECT 2191.630 3098.590 2192.810 3099.770 ;
        RECT 2193.230 3098.590 2194.410 3099.770 ;
        RECT 2191.630 3096.990 2192.810 3098.170 ;
        RECT 2193.230 3096.990 2194.410 3098.170 ;
        RECT 2191.630 2918.590 2192.810 2919.770 ;
        RECT 2193.230 2918.590 2194.410 2919.770 ;
        RECT 2191.630 2916.990 2192.810 2918.170 ;
        RECT 2193.230 2916.990 2194.410 2918.170 ;
        RECT 2191.630 2738.590 2192.810 2739.770 ;
        RECT 2193.230 2738.590 2194.410 2739.770 ;
        RECT 2191.630 2736.990 2192.810 2738.170 ;
        RECT 2193.230 2736.990 2194.410 2738.170 ;
        RECT 2191.630 2558.590 2192.810 2559.770 ;
        RECT 2193.230 2558.590 2194.410 2559.770 ;
        RECT 2191.630 2556.990 2192.810 2558.170 ;
        RECT 2193.230 2556.990 2194.410 2558.170 ;
        RECT 2191.630 2378.590 2192.810 2379.770 ;
        RECT 2193.230 2378.590 2194.410 2379.770 ;
        RECT 2191.630 2376.990 2192.810 2378.170 ;
        RECT 2193.230 2376.990 2194.410 2378.170 ;
        RECT 2191.630 2198.590 2192.810 2199.770 ;
        RECT 2193.230 2198.590 2194.410 2199.770 ;
        RECT 2191.630 2196.990 2192.810 2198.170 ;
        RECT 2193.230 2196.990 2194.410 2198.170 ;
        RECT 2191.630 2018.590 2192.810 2019.770 ;
        RECT 2193.230 2018.590 2194.410 2019.770 ;
        RECT 2191.630 2016.990 2192.810 2018.170 ;
        RECT 2193.230 2016.990 2194.410 2018.170 ;
        RECT 2191.630 1838.590 2192.810 1839.770 ;
        RECT 2193.230 1838.590 2194.410 1839.770 ;
        RECT 2191.630 1836.990 2192.810 1838.170 ;
        RECT 2193.230 1836.990 2194.410 1838.170 ;
        RECT 2191.630 1658.590 2192.810 1659.770 ;
        RECT 2193.230 1658.590 2194.410 1659.770 ;
        RECT 2191.630 1656.990 2192.810 1658.170 ;
        RECT 2193.230 1656.990 2194.410 1658.170 ;
        RECT 2191.630 1478.590 2192.810 1479.770 ;
        RECT 2193.230 1478.590 2194.410 1479.770 ;
        RECT 2191.630 1476.990 2192.810 1478.170 ;
        RECT 2193.230 1476.990 2194.410 1478.170 ;
        RECT 2191.630 1298.590 2192.810 1299.770 ;
        RECT 2193.230 1298.590 2194.410 1299.770 ;
        RECT 2191.630 1296.990 2192.810 1298.170 ;
        RECT 2193.230 1296.990 2194.410 1298.170 ;
        RECT 2191.630 1118.590 2192.810 1119.770 ;
        RECT 2193.230 1118.590 2194.410 1119.770 ;
        RECT 2191.630 1116.990 2192.810 1118.170 ;
        RECT 2193.230 1116.990 2194.410 1118.170 ;
        RECT 2191.630 938.590 2192.810 939.770 ;
        RECT 2193.230 938.590 2194.410 939.770 ;
        RECT 2191.630 936.990 2192.810 938.170 ;
        RECT 2193.230 936.990 2194.410 938.170 ;
        RECT 2191.630 758.590 2192.810 759.770 ;
        RECT 2193.230 758.590 2194.410 759.770 ;
        RECT 2191.630 756.990 2192.810 758.170 ;
        RECT 2193.230 756.990 2194.410 758.170 ;
        RECT 2191.630 578.590 2192.810 579.770 ;
        RECT 2193.230 578.590 2194.410 579.770 ;
        RECT 2191.630 576.990 2192.810 578.170 ;
        RECT 2193.230 576.990 2194.410 578.170 ;
        RECT 2191.630 398.590 2192.810 399.770 ;
        RECT 2193.230 398.590 2194.410 399.770 ;
        RECT 2191.630 396.990 2192.810 398.170 ;
        RECT 2193.230 396.990 2194.410 398.170 ;
        RECT 2191.630 218.590 2192.810 219.770 ;
        RECT 2193.230 218.590 2194.410 219.770 ;
        RECT 2191.630 216.990 2192.810 218.170 ;
        RECT 2193.230 216.990 2194.410 218.170 ;
        RECT 2191.630 38.590 2192.810 39.770 ;
        RECT 2193.230 38.590 2194.410 39.770 ;
        RECT 2191.630 36.990 2192.810 38.170 ;
        RECT 2193.230 36.990 2194.410 38.170 ;
        RECT 2191.630 -7.710 2192.810 -6.530 ;
        RECT 2193.230 -7.710 2194.410 -6.530 ;
        RECT 2191.630 -9.310 2192.810 -8.130 ;
        RECT 2193.230 -9.310 2194.410 -8.130 ;
        RECT 2371.630 3527.810 2372.810 3528.990 ;
        RECT 2373.230 3527.810 2374.410 3528.990 ;
        RECT 2371.630 3526.210 2372.810 3527.390 ;
        RECT 2373.230 3526.210 2374.410 3527.390 ;
        RECT 2371.630 3458.590 2372.810 3459.770 ;
        RECT 2373.230 3458.590 2374.410 3459.770 ;
        RECT 2371.630 3456.990 2372.810 3458.170 ;
        RECT 2373.230 3456.990 2374.410 3458.170 ;
        RECT 2371.630 3278.590 2372.810 3279.770 ;
        RECT 2373.230 3278.590 2374.410 3279.770 ;
        RECT 2371.630 3276.990 2372.810 3278.170 ;
        RECT 2373.230 3276.990 2374.410 3278.170 ;
        RECT 2371.630 3098.590 2372.810 3099.770 ;
        RECT 2373.230 3098.590 2374.410 3099.770 ;
        RECT 2371.630 3096.990 2372.810 3098.170 ;
        RECT 2373.230 3096.990 2374.410 3098.170 ;
        RECT 2371.630 2918.590 2372.810 2919.770 ;
        RECT 2373.230 2918.590 2374.410 2919.770 ;
        RECT 2371.630 2916.990 2372.810 2918.170 ;
        RECT 2373.230 2916.990 2374.410 2918.170 ;
        RECT 2371.630 2738.590 2372.810 2739.770 ;
        RECT 2373.230 2738.590 2374.410 2739.770 ;
        RECT 2371.630 2736.990 2372.810 2738.170 ;
        RECT 2373.230 2736.990 2374.410 2738.170 ;
        RECT 2371.630 2558.590 2372.810 2559.770 ;
        RECT 2373.230 2558.590 2374.410 2559.770 ;
        RECT 2371.630 2556.990 2372.810 2558.170 ;
        RECT 2373.230 2556.990 2374.410 2558.170 ;
        RECT 2371.630 2378.590 2372.810 2379.770 ;
        RECT 2373.230 2378.590 2374.410 2379.770 ;
        RECT 2371.630 2376.990 2372.810 2378.170 ;
        RECT 2373.230 2376.990 2374.410 2378.170 ;
        RECT 2371.630 2198.590 2372.810 2199.770 ;
        RECT 2373.230 2198.590 2374.410 2199.770 ;
        RECT 2371.630 2196.990 2372.810 2198.170 ;
        RECT 2373.230 2196.990 2374.410 2198.170 ;
        RECT 2371.630 2018.590 2372.810 2019.770 ;
        RECT 2373.230 2018.590 2374.410 2019.770 ;
        RECT 2371.630 2016.990 2372.810 2018.170 ;
        RECT 2373.230 2016.990 2374.410 2018.170 ;
        RECT 2371.630 1838.590 2372.810 1839.770 ;
        RECT 2373.230 1838.590 2374.410 1839.770 ;
        RECT 2371.630 1836.990 2372.810 1838.170 ;
        RECT 2373.230 1836.990 2374.410 1838.170 ;
        RECT 2371.630 1658.590 2372.810 1659.770 ;
        RECT 2373.230 1658.590 2374.410 1659.770 ;
        RECT 2371.630 1656.990 2372.810 1658.170 ;
        RECT 2373.230 1656.990 2374.410 1658.170 ;
        RECT 2371.630 1478.590 2372.810 1479.770 ;
        RECT 2373.230 1478.590 2374.410 1479.770 ;
        RECT 2371.630 1476.990 2372.810 1478.170 ;
        RECT 2373.230 1476.990 2374.410 1478.170 ;
        RECT 2371.630 1298.590 2372.810 1299.770 ;
        RECT 2373.230 1298.590 2374.410 1299.770 ;
        RECT 2371.630 1296.990 2372.810 1298.170 ;
        RECT 2373.230 1296.990 2374.410 1298.170 ;
        RECT 2371.630 1118.590 2372.810 1119.770 ;
        RECT 2373.230 1118.590 2374.410 1119.770 ;
        RECT 2371.630 1116.990 2372.810 1118.170 ;
        RECT 2373.230 1116.990 2374.410 1118.170 ;
        RECT 2371.630 938.590 2372.810 939.770 ;
        RECT 2373.230 938.590 2374.410 939.770 ;
        RECT 2371.630 936.990 2372.810 938.170 ;
        RECT 2373.230 936.990 2374.410 938.170 ;
        RECT 2371.630 758.590 2372.810 759.770 ;
        RECT 2373.230 758.590 2374.410 759.770 ;
        RECT 2371.630 756.990 2372.810 758.170 ;
        RECT 2373.230 756.990 2374.410 758.170 ;
        RECT 2371.630 578.590 2372.810 579.770 ;
        RECT 2373.230 578.590 2374.410 579.770 ;
        RECT 2371.630 576.990 2372.810 578.170 ;
        RECT 2373.230 576.990 2374.410 578.170 ;
        RECT 2371.630 398.590 2372.810 399.770 ;
        RECT 2373.230 398.590 2374.410 399.770 ;
        RECT 2371.630 396.990 2372.810 398.170 ;
        RECT 2373.230 396.990 2374.410 398.170 ;
        RECT 2371.630 218.590 2372.810 219.770 ;
        RECT 2373.230 218.590 2374.410 219.770 ;
        RECT 2371.630 216.990 2372.810 218.170 ;
        RECT 2373.230 216.990 2374.410 218.170 ;
        RECT 2371.630 38.590 2372.810 39.770 ;
        RECT 2373.230 38.590 2374.410 39.770 ;
        RECT 2371.630 36.990 2372.810 38.170 ;
        RECT 2373.230 36.990 2374.410 38.170 ;
        RECT 2371.630 -7.710 2372.810 -6.530 ;
        RECT 2373.230 -7.710 2374.410 -6.530 ;
        RECT 2371.630 -9.310 2372.810 -8.130 ;
        RECT 2373.230 -9.310 2374.410 -8.130 ;
        RECT 2551.630 3527.810 2552.810 3528.990 ;
        RECT 2553.230 3527.810 2554.410 3528.990 ;
        RECT 2551.630 3526.210 2552.810 3527.390 ;
        RECT 2553.230 3526.210 2554.410 3527.390 ;
        RECT 2551.630 3458.590 2552.810 3459.770 ;
        RECT 2553.230 3458.590 2554.410 3459.770 ;
        RECT 2551.630 3456.990 2552.810 3458.170 ;
        RECT 2553.230 3456.990 2554.410 3458.170 ;
        RECT 2551.630 3278.590 2552.810 3279.770 ;
        RECT 2553.230 3278.590 2554.410 3279.770 ;
        RECT 2551.630 3276.990 2552.810 3278.170 ;
        RECT 2553.230 3276.990 2554.410 3278.170 ;
        RECT 2551.630 3098.590 2552.810 3099.770 ;
        RECT 2553.230 3098.590 2554.410 3099.770 ;
        RECT 2551.630 3096.990 2552.810 3098.170 ;
        RECT 2553.230 3096.990 2554.410 3098.170 ;
        RECT 2551.630 2918.590 2552.810 2919.770 ;
        RECT 2553.230 2918.590 2554.410 2919.770 ;
        RECT 2551.630 2916.990 2552.810 2918.170 ;
        RECT 2553.230 2916.990 2554.410 2918.170 ;
        RECT 2551.630 2738.590 2552.810 2739.770 ;
        RECT 2553.230 2738.590 2554.410 2739.770 ;
        RECT 2551.630 2736.990 2552.810 2738.170 ;
        RECT 2553.230 2736.990 2554.410 2738.170 ;
        RECT 2551.630 2558.590 2552.810 2559.770 ;
        RECT 2553.230 2558.590 2554.410 2559.770 ;
        RECT 2551.630 2556.990 2552.810 2558.170 ;
        RECT 2553.230 2556.990 2554.410 2558.170 ;
        RECT 2551.630 2378.590 2552.810 2379.770 ;
        RECT 2553.230 2378.590 2554.410 2379.770 ;
        RECT 2551.630 2376.990 2552.810 2378.170 ;
        RECT 2553.230 2376.990 2554.410 2378.170 ;
        RECT 2551.630 2198.590 2552.810 2199.770 ;
        RECT 2553.230 2198.590 2554.410 2199.770 ;
        RECT 2551.630 2196.990 2552.810 2198.170 ;
        RECT 2553.230 2196.990 2554.410 2198.170 ;
        RECT 2551.630 2018.590 2552.810 2019.770 ;
        RECT 2553.230 2018.590 2554.410 2019.770 ;
        RECT 2551.630 2016.990 2552.810 2018.170 ;
        RECT 2553.230 2016.990 2554.410 2018.170 ;
        RECT 2551.630 1838.590 2552.810 1839.770 ;
        RECT 2553.230 1838.590 2554.410 1839.770 ;
        RECT 2551.630 1836.990 2552.810 1838.170 ;
        RECT 2553.230 1836.990 2554.410 1838.170 ;
        RECT 2551.630 1658.590 2552.810 1659.770 ;
        RECT 2553.230 1658.590 2554.410 1659.770 ;
        RECT 2551.630 1656.990 2552.810 1658.170 ;
        RECT 2553.230 1656.990 2554.410 1658.170 ;
        RECT 2551.630 1478.590 2552.810 1479.770 ;
        RECT 2553.230 1478.590 2554.410 1479.770 ;
        RECT 2551.630 1476.990 2552.810 1478.170 ;
        RECT 2553.230 1476.990 2554.410 1478.170 ;
        RECT 2551.630 1298.590 2552.810 1299.770 ;
        RECT 2553.230 1298.590 2554.410 1299.770 ;
        RECT 2551.630 1296.990 2552.810 1298.170 ;
        RECT 2553.230 1296.990 2554.410 1298.170 ;
        RECT 2551.630 1118.590 2552.810 1119.770 ;
        RECT 2553.230 1118.590 2554.410 1119.770 ;
        RECT 2551.630 1116.990 2552.810 1118.170 ;
        RECT 2553.230 1116.990 2554.410 1118.170 ;
        RECT 2551.630 938.590 2552.810 939.770 ;
        RECT 2553.230 938.590 2554.410 939.770 ;
        RECT 2551.630 936.990 2552.810 938.170 ;
        RECT 2553.230 936.990 2554.410 938.170 ;
        RECT 2551.630 758.590 2552.810 759.770 ;
        RECT 2553.230 758.590 2554.410 759.770 ;
        RECT 2551.630 756.990 2552.810 758.170 ;
        RECT 2553.230 756.990 2554.410 758.170 ;
        RECT 2551.630 578.590 2552.810 579.770 ;
        RECT 2553.230 578.590 2554.410 579.770 ;
        RECT 2551.630 576.990 2552.810 578.170 ;
        RECT 2553.230 576.990 2554.410 578.170 ;
        RECT 2551.630 398.590 2552.810 399.770 ;
        RECT 2553.230 398.590 2554.410 399.770 ;
        RECT 2551.630 396.990 2552.810 398.170 ;
        RECT 2553.230 396.990 2554.410 398.170 ;
        RECT 2551.630 218.590 2552.810 219.770 ;
        RECT 2553.230 218.590 2554.410 219.770 ;
        RECT 2551.630 216.990 2552.810 218.170 ;
        RECT 2553.230 216.990 2554.410 218.170 ;
        RECT 2551.630 38.590 2552.810 39.770 ;
        RECT 2553.230 38.590 2554.410 39.770 ;
        RECT 2551.630 36.990 2552.810 38.170 ;
        RECT 2553.230 36.990 2554.410 38.170 ;
        RECT 2551.630 -7.710 2552.810 -6.530 ;
        RECT 2553.230 -7.710 2554.410 -6.530 ;
        RECT 2551.630 -9.310 2552.810 -8.130 ;
        RECT 2553.230 -9.310 2554.410 -8.130 ;
        RECT 2731.630 3527.810 2732.810 3528.990 ;
        RECT 2733.230 3527.810 2734.410 3528.990 ;
        RECT 2731.630 3526.210 2732.810 3527.390 ;
        RECT 2733.230 3526.210 2734.410 3527.390 ;
        RECT 2731.630 3458.590 2732.810 3459.770 ;
        RECT 2733.230 3458.590 2734.410 3459.770 ;
        RECT 2731.630 3456.990 2732.810 3458.170 ;
        RECT 2733.230 3456.990 2734.410 3458.170 ;
        RECT 2731.630 3278.590 2732.810 3279.770 ;
        RECT 2733.230 3278.590 2734.410 3279.770 ;
        RECT 2731.630 3276.990 2732.810 3278.170 ;
        RECT 2733.230 3276.990 2734.410 3278.170 ;
        RECT 2731.630 3098.590 2732.810 3099.770 ;
        RECT 2733.230 3098.590 2734.410 3099.770 ;
        RECT 2731.630 3096.990 2732.810 3098.170 ;
        RECT 2733.230 3096.990 2734.410 3098.170 ;
        RECT 2731.630 2918.590 2732.810 2919.770 ;
        RECT 2733.230 2918.590 2734.410 2919.770 ;
        RECT 2731.630 2916.990 2732.810 2918.170 ;
        RECT 2733.230 2916.990 2734.410 2918.170 ;
        RECT 2731.630 2738.590 2732.810 2739.770 ;
        RECT 2733.230 2738.590 2734.410 2739.770 ;
        RECT 2731.630 2736.990 2732.810 2738.170 ;
        RECT 2733.230 2736.990 2734.410 2738.170 ;
        RECT 2731.630 2558.590 2732.810 2559.770 ;
        RECT 2733.230 2558.590 2734.410 2559.770 ;
        RECT 2731.630 2556.990 2732.810 2558.170 ;
        RECT 2733.230 2556.990 2734.410 2558.170 ;
        RECT 2731.630 2378.590 2732.810 2379.770 ;
        RECT 2733.230 2378.590 2734.410 2379.770 ;
        RECT 2731.630 2376.990 2732.810 2378.170 ;
        RECT 2733.230 2376.990 2734.410 2378.170 ;
        RECT 2731.630 2198.590 2732.810 2199.770 ;
        RECT 2733.230 2198.590 2734.410 2199.770 ;
        RECT 2731.630 2196.990 2732.810 2198.170 ;
        RECT 2733.230 2196.990 2734.410 2198.170 ;
        RECT 2731.630 2018.590 2732.810 2019.770 ;
        RECT 2733.230 2018.590 2734.410 2019.770 ;
        RECT 2731.630 2016.990 2732.810 2018.170 ;
        RECT 2733.230 2016.990 2734.410 2018.170 ;
        RECT 2731.630 1838.590 2732.810 1839.770 ;
        RECT 2733.230 1838.590 2734.410 1839.770 ;
        RECT 2731.630 1836.990 2732.810 1838.170 ;
        RECT 2733.230 1836.990 2734.410 1838.170 ;
        RECT 2731.630 1658.590 2732.810 1659.770 ;
        RECT 2733.230 1658.590 2734.410 1659.770 ;
        RECT 2731.630 1656.990 2732.810 1658.170 ;
        RECT 2733.230 1656.990 2734.410 1658.170 ;
        RECT 2731.630 1478.590 2732.810 1479.770 ;
        RECT 2733.230 1478.590 2734.410 1479.770 ;
        RECT 2731.630 1476.990 2732.810 1478.170 ;
        RECT 2733.230 1476.990 2734.410 1478.170 ;
        RECT 2731.630 1298.590 2732.810 1299.770 ;
        RECT 2733.230 1298.590 2734.410 1299.770 ;
        RECT 2731.630 1296.990 2732.810 1298.170 ;
        RECT 2733.230 1296.990 2734.410 1298.170 ;
        RECT 2731.630 1118.590 2732.810 1119.770 ;
        RECT 2733.230 1118.590 2734.410 1119.770 ;
        RECT 2731.630 1116.990 2732.810 1118.170 ;
        RECT 2733.230 1116.990 2734.410 1118.170 ;
        RECT 2731.630 938.590 2732.810 939.770 ;
        RECT 2733.230 938.590 2734.410 939.770 ;
        RECT 2731.630 936.990 2732.810 938.170 ;
        RECT 2733.230 936.990 2734.410 938.170 ;
        RECT 2731.630 758.590 2732.810 759.770 ;
        RECT 2733.230 758.590 2734.410 759.770 ;
        RECT 2731.630 756.990 2732.810 758.170 ;
        RECT 2733.230 756.990 2734.410 758.170 ;
        RECT 2731.630 578.590 2732.810 579.770 ;
        RECT 2733.230 578.590 2734.410 579.770 ;
        RECT 2731.630 576.990 2732.810 578.170 ;
        RECT 2733.230 576.990 2734.410 578.170 ;
        RECT 2731.630 398.590 2732.810 399.770 ;
        RECT 2733.230 398.590 2734.410 399.770 ;
        RECT 2731.630 396.990 2732.810 398.170 ;
        RECT 2733.230 396.990 2734.410 398.170 ;
        RECT 2731.630 218.590 2732.810 219.770 ;
        RECT 2733.230 218.590 2734.410 219.770 ;
        RECT 2731.630 216.990 2732.810 218.170 ;
        RECT 2733.230 216.990 2734.410 218.170 ;
        RECT 2731.630 38.590 2732.810 39.770 ;
        RECT 2733.230 38.590 2734.410 39.770 ;
        RECT 2731.630 36.990 2732.810 38.170 ;
        RECT 2733.230 36.990 2734.410 38.170 ;
        RECT 2731.630 -7.710 2732.810 -6.530 ;
        RECT 2733.230 -7.710 2734.410 -6.530 ;
        RECT 2731.630 -9.310 2732.810 -8.130 ;
        RECT 2733.230 -9.310 2734.410 -8.130 ;
        RECT 2911.630 3527.810 2912.810 3528.990 ;
        RECT 2913.230 3527.810 2914.410 3528.990 ;
        RECT 2911.630 3526.210 2912.810 3527.390 ;
        RECT 2913.230 3526.210 2914.410 3527.390 ;
        RECT 2911.630 3458.590 2912.810 3459.770 ;
        RECT 2913.230 3458.590 2914.410 3459.770 ;
        RECT 2911.630 3456.990 2912.810 3458.170 ;
        RECT 2913.230 3456.990 2914.410 3458.170 ;
        RECT 2911.630 3278.590 2912.810 3279.770 ;
        RECT 2913.230 3278.590 2914.410 3279.770 ;
        RECT 2911.630 3276.990 2912.810 3278.170 ;
        RECT 2913.230 3276.990 2914.410 3278.170 ;
        RECT 2911.630 3098.590 2912.810 3099.770 ;
        RECT 2913.230 3098.590 2914.410 3099.770 ;
        RECT 2911.630 3096.990 2912.810 3098.170 ;
        RECT 2913.230 3096.990 2914.410 3098.170 ;
        RECT 2911.630 2918.590 2912.810 2919.770 ;
        RECT 2913.230 2918.590 2914.410 2919.770 ;
        RECT 2911.630 2916.990 2912.810 2918.170 ;
        RECT 2913.230 2916.990 2914.410 2918.170 ;
        RECT 2911.630 2738.590 2912.810 2739.770 ;
        RECT 2913.230 2738.590 2914.410 2739.770 ;
        RECT 2911.630 2736.990 2912.810 2738.170 ;
        RECT 2913.230 2736.990 2914.410 2738.170 ;
        RECT 2911.630 2558.590 2912.810 2559.770 ;
        RECT 2913.230 2558.590 2914.410 2559.770 ;
        RECT 2911.630 2556.990 2912.810 2558.170 ;
        RECT 2913.230 2556.990 2914.410 2558.170 ;
        RECT 2911.630 2378.590 2912.810 2379.770 ;
        RECT 2913.230 2378.590 2914.410 2379.770 ;
        RECT 2911.630 2376.990 2912.810 2378.170 ;
        RECT 2913.230 2376.990 2914.410 2378.170 ;
        RECT 2911.630 2198.590 2912.810 2199.770 ;
        RECT 2913.230 2198.590 2914.410 2199.770 ;
        RECT 2911.630 2196.990 2912.810 2198.170 ;
        RECT 2913.230 2196.990 2914.410 2198.170 ;
        RECT 2911.630 2018.590 2912.810 2019.770 ;
        RECT 2913.230 2018.590 2914.410 2019.770 ;
        RECT 2911.630 2016.990 2912.810 2018.170 ;
        RECT 2913.230 2016.990 2914.410 2018.170 ;
        RECT 2911.630 1838.590 2912.810 1839.770 ;
        RECT 2913.230 1838.590 2914.410 1839.770 ;
        RECT 2911.630 1836.990 2912.810 1838.170 ;
        RECT 2913.230 1836.990 2914.410 1838.170 ;
        RECT 2911.630 1658.590 2912.810 1659.770 ;
        RECT 2913.230 1658.590 2914.410 1659.770 ;
        RECT 2911.630 1656.990 2912.810 1658.170 ;
        RECT 2913.230 1656.990 2914.410 1658.170 ;
        RECT 2911.630 1478.590 2912.810 1479.770 ;
        RECT 2913.230 1478.590 2914.410 1479.770 ;
        RECT 2911.630 1476.990 2912.810 1478.170 ;
        RECT 2913.230 1476.990 2914.410 1478.170 ;
        RECT 2911.630 1298.590 2912.810 1299.770 ;
        RECT 2913.230 1298.590 2914.410 1299.770 ;
        RECT 2911.630 1296.990 2912.810 1298.170 ;
        RECT 2913.230 1296.990 2914.410 1298.170 ;
        RECT 2911.630 1118.590 2912.810 1119.770 ;
        RECT 2913.230 1118.590 2914.410 1119.770 ;
        RECT 2911.630 1116.990 2912.810 1118.170 ;
        RECT 2913.230 1116.990 2914.410 1118.170 ;
        RECT 2911.630 938.590 2912.810 939.770 ;
        RECT 2913.230 938.590 2914.410 939.770 ;
        RECT 2911.630 936.990 2912.810 938.170 ;
        RECT 2913.230 936.990 2914.410 938.170 ;
        RECT 2911.630 758.590 2912.810 759.770 ;
        RECT 2913.230 758.590 2914.410 759.770 ;
        RECT 2911.630 756.990 2912.810 758.170 ;
        RECT 2913.230 756.990 2914.410 758.170 ;
        RECT 2911.630 578.590 2912.810 579.770 ;
        RECT 2913.230 578.590 2914.410 579.770 ;
        RECT 2911.630 576.990 2912.810 578.170 ;
        RECT 2913.230 576.990 2914.410 578.170 ;
        RECT 2911.630 398.590 2912.810 399.770 ;
        RECT 2913.230 398.590 2914.410 399.770 ;
        RECT 2911.630 396.990 2912.810 398.170 ;
        RECT 2913.230 396.990 2914.410 398.170 ;
        RECT 2911.630 218.590 2912.810 219.770 ;
        RECT 2913.230 218.590 2914.410 219.770 ;
        RECT 2911.630 216.990 2912.810 218.170 ;
        RECT 2913.230 216.990 2914.410 218.170 ;
        RECT 2911.630 38.590 2912.810 39.770 ;
        RECT 2913.230 38.590 2914.410 39.770 ;
        RECT 2911.630 36.990 2912.810 38.170 ;
        RECT 2913.230 36.990 2914.410 38.170 ;
        RECT 2911.630 -7.710 2912.810 -6.530 ;
        RECT 2913.230 -7.710 2914.410 -6.530 ;
        RECT 2911.630 -9.310 2912.810 -8.130 ;
        RECT 2913.230 -9.310 2914.410 -8.130 ;
        RECT 2931.510 3527.810 2932.690 3528.990 ;
        RECT 2933.110 3527.810 2934.290 3528.990 ;
        RECT 2931.510 3526.210 2932.690 3527.390 ;
        RECT 2933.110 3526.210 2934.290 3527.390 ;
        RECT 2931.510 3458.590 2932.690 3459.770 ;
        RECT 2933.110 3458.590 2934.290 3459.770 ;
        RECT 2931.510 3456.990 2932.690 3458.170 ;
        RECT 2933.110 3456.990 2934.290 3458.170 ;
        RECT 2931.510 3278.590 2932.690 3279.770 ;
        RECT 2933.110 3278.590 2934.290 3279.770 ;
        RECT 2931.510 3276.990 2932.690 3278.170 ;
        RECT 2933.110 3276.990 2934.290 3278.170 ;
        RECT 2931.510 3098.590 2932.690 3099.770 ;
        RECT 2933.110 3098.590 2934.290 3099.770 ;
        RECT 2931.510 3096.990 2932.690 3098.170 ;
        RECT 2933.110 3096.990 2934.290 3098.170 ;
        RECT 2931.510 2918.590 2932.690 2919.770 ;
        RECT 2933.110 2918.590 2934.290 2919.770 ;
        RECT 2931.510 2916.990 2932.690 2918.170 ;
        RECT 2933.110 2916.990 2934.290 2918.170 ;
        RECT 2931.510 2738.590 2932.690 2739.770 ;
        RECT 2933.110 2738.590 2934.290 2739.770 ;
        RECT 2931.510 2736.990 2932.690 2738.170 ;
        RECT 2933.110 2736.990 2934.290 2738.170 ;
        RECT 2931.510 2558.590 2932.690 2559.770 ;
        RECT 2933.110 2558.590 2934.290 2559.770 ;
        RECT 2931.510 2556.990 2932.690 2558.170 ;
        RECT 2933.110 2556.990 2934.290 2558.170 ;
        RECT 2931.510 2378.590 2932.690 2379.770 ;
        RECT 2933.110 2378.590 2934.290 2379.770 ;
        RECT 2931.510 2376.990 2932.690 2378.170 ;
        RECT 2933.110 2376.990 2934.290 2378.170 ;
        RECT 2931.510 2198.590 2932.690 2199.770 ;
        RECT 2933.110 2198.590 2934.290 2199.770 ;
        RECT 2931.510 2196.990 2932.690 2198.170 ;
        RECT 2933.110 2196.990 2934.290 2198.170 ;
        RECT 2931.510 2018.590 2932.690 2019.770 ;
        RECT 2933.110 2018.590 2934.290 2019.770 ;
        RECT 2931.510 2016.990 2932.690 2018.170 ;
        RECT 2933.110 2016.990 2934.290 2018.170 ;
        RECT 2931.510 1838.590 2932.690 1839.770 ;
        RECT 2933.110 1838.590 2934.290 1839.770 ;
        RECT 2931.510 1836.990 2932.690 1838.170 ;
        RECT 2933.110 1836.990 2934.290 1838.170 ;
        RECT 2931.510 1658.590 2932.690 1659.770 ;
        RECT 2933.110 1658.590 2934.290 1659.770 ;
        RECT 2931.510 1656.990 2932.690 1658.170 ;
        RECT 2933.110 1656.990 2934.290 1658.170 ;
        RECT 2931.510 1478.590 2932.690 1479.770 ;
        RECT 2933.110 1478.590 2934.290 1479.770 ;
        RECT 2931.510 1476.990 2932.690 1478.170 ;
        RECT 2933.110 1476.990 2934.290 1478.170 ;
        RECT 2931.510 1298.590 2932.690 1299.770 ;
        RECT 2933.110 1298.590 2934.290 1299.770 ;
        RECT 2931.510 1296.990 2932.690 1298.170 ;
        RECT 2933.110 1296.990 2934.290 1298.170 ;
        RECT 2931.510 1118.590 2932.690 1119.770 ;
        RECT 2933.110 1118.590 2934.290 1119.770 ;
        RECT 2931.510 1116.990 2932.690 1118.170 ;
        RECT 2933.110 1116.990 2934.290 1118.170 ;
        RECT 2931.510 938.590 2932.690 939.770 ;
        RECT 2933.110 938.590 2934.290 939.770 ;
        RECT 2931.510 936.990 2932.690 938.170 ;
        RECT 2933.110 936.990 2934.290 938.170 ;
        RECT 2931.510 758.590 2932.690 759.770 ;
        RECT 2933.110 758.590 2934.290 759.770 ;
        RECT 2931.510 756.990 2932.690 758.170 ;
        RECT 2933.110 756.990 2934.290 758.170 ;
        RECT 2931.510 578.590 2932.690 579.770 ;
        RECT 2933.110 578.590 2934.290 579.770 ;
        RECT 2931.510 576.990 2932.690 578.170 ;
        RECT 2933.110 576.990 2934.290 578.170 ;
        RECT 2931.510 398.590 2932.690 399.770 ;
        RECT 2933.110 398.590 2934.290 399.770 ;
        RECT 2931.510 396.990 2932.690 398.170 ;
        RECT 2933.110 396.990 2934.290 398.170 ;
        RECT 2931.510 218.590 2932.690 219.770 ;
        RECT 2933.110 218.590 2934.290 219.770 ;
        RECT 2931.510 216.990 2932.690 218.170 ;
        RECT 2933.110 216.990 2934.290 218.170 ;
        RECT 2931.510 38.590 2932.690 39.770 ;
        RECT 2933.110 38.590 2934.290 39.770 ;
        RECT 2931.510 36.990 2932.690 38.170 ;
        RECT 2933.110 36.990 2934.290 38.170 ;
        RECT 2931.510 -7.710 2932.690 -6.530 ;
        RECT 2933.110 -7.710 2934.290 -6.530 ;
        RECT 2931.510 -9.310 2932.690 -8.130 ;
        RECT 2933.110 -9.310 2934.290 -8.130 ;
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
        RECT -43.630 3456.830 2963.250 3459.930 ;
        RECT -43.630 3276.830 2963.250 3279.930 ;
        RECT -43.630 3096.830 2963.250 3099.930 ;
        RECT -43.630 2916.830 2963.250 2919.930 ;
        RECT -43.630 2736.830 2963.250 2739.930 ;
        RECT -43.630 2556.830 2963.250 2559.930 ;
        RECT -43.630 2376.830 2963.250 2379.930 ;
        RECT -43.630 2196.830 2963.250 2199.930 ;
        RECT -43.630 2016.830 2963.250 2019.930 ;
        RECT -43.630 1836.830 2963.250 1839.930 ;
        RECT -43.630 1656.830 2963.250 1659.930 ;
        RECT -43.630 1476.830 2963.250 1479.930 ;
        RECT -43.630 1296.830 2963.250 1299.930 ;
        RECT -43.630 1116.830 2963.250 1119.930 ;
        RECT -43.630 936.830 2963.250 939.930 ;
        RECT -43.630 756.830 2963.250 759.930 ;
        RECT -43.630 576.830 2963.250 579.930 ;
        RECT -43.630 396.830 2963.250 399.930 ;
        RECT -43.630 216.830 2963.250 219.930 ;
        RECT -43.630 36.830 2963.250 39.930 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
        RECT 76.470 -38.270 79.570 3557.950 ;
        RECT 256.470 -38.270 259.570 3557.950 ;
        RECT 436.470 810.000 439.570 3557.950 ;
        RECT 616.470 810.000 619.570 3557.950 ;
        RECT 436.470 -38.270 439.570 490.000 ;
        RECT 616.470 -38.270 619.570 490.000 ;
        RECT 796.470 -38.270 799.570 3557.950 ;
        RECT 976.470 -38.270 979.570 3557.950 ;
        RECT 1156.470 -38.270 1159.570 3557.950 ;
        RECT 1336.470 -38.270 1339.570 3557.950 ;
        RECT 1516.470 -38.270 1519.570 3557.950 ;
        RECT 1696.470 -38.270 1699.570 3557.950 ;
        RECT 1876.470 -38.270 1879.570 3557.950 ;
        RECT 2056.470 -38.270 2059.570 3557.950 ;
        RECT 2236.470 -38.270 2239.570 3557.950 ;
        RECT 2416.470 -38.270 2419.570 3557.950 ;
        RECT 2596.470 -38.270 2599.570 3557.950 ;
        RECT 2776.470 -38.270 2779.570 3557.950 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
      LAYER via4 ;
        RECT -24.270 3537.410 -23.090 3538.590 ;
        RECT -22.670 3537.410 -21.490 3538.590 ;
        RECT -24.270 3535.810 -23.090 3536.990 ;
        RECT -22.670 3535.810 -21.490 3536.990 ;
        RECT -24.270 3503.590 -23.090 3504.770 ;
        RECT -22.670 3503.590 -21.490 3504.770 ;
        RECT -24.270 3501.990 -23.090 3503.170 ;
        RECT -22.670 3501.990 -21.490 3503.170 ;
        RECT -24.270 3323.590 -23.090 3324.770 ;
        RECT -22.670 3323.590 -21.490 3324.770 ;
        RECT -24.270 3321.990 -23.090 3323.170 ;
        RECT -22.670 3321.990 -21.490 3323.170 ;
        RECT -24.270 3143.590 -23.090 3144.770 ;
        RECT -22.670 3143.590 -21.490 3144.770 ;
        RECT -24.270 3141.990 -23.090 3143.170 ;
        RECT -22.670 3141.990 -21.490 3143.170 ;
        RECT -24.270 2963.590 -23.090 2964.770 ;
        RECT -22.670 2963.590 -21.490 2964.770 ;
        RECT -24.270 2961.990 -23.090 2963.170 ;
        RECT -22.670 2961.990 -21.490 2963.170 ;
        RECT -24.270 2783.590 -23.090 2784.770 ;
        RECT -22.670 2783.590 -21.490 2784.770 ;
        RECT -24.270 2781.990 -23.090 2783.170 ;
        RECT -22.670 2781.990 -21.490 2783.170 ;
        RECT -24.270 2603.590 -23.090 2604.770 ;
        RECT -22.670 2603.590 -21.490 2604.770 ;
        RECT -24.270 2601.990 -23.090 2603.170 ;
        RECT -22.670 2601.990 -21.490 2603.170 ;
        RECT -24.270 2423.590 -23.090 2424.770 ;
        RECT -22.670 2423.590 -21.490 2424.770 ;
        RECT -24.270 2421.990 -23.090 2423.170 ;
        RECT -22.670 2421.990 -21.490 2423.170 ;
        RECT -24.270 2243.590 -23.090 2244.770 ;
        RECT -22.670 2243.590 -21.490 2244.770 ;
        RECT -24.270 2241.990 -23.090 2243.170 ;
        RECT -22.670 2241.990 -21.490 2243.170 ;
        RECT -24.270 2063.590 -23.090 2064.770 ;
        RECT -22.670 2063.590 -21.490 2064.770 ;
        RECT -24.270 2061.990 -23.090 2063.170 ;
        RECT -22.670 2061.990 -21.490 2063.170 ;
        RECT -24.270 1883.590 -23.090 1884.770 ;
        RECT -22.670 1883.590 -21.490 1884.770 ;
        RECT -24.270 1881.990 -23.090 1883.170 ;
        RECT -22.670 1881.990 -21.490 1883.170 ;
        RECT -24.270 1703.590 -23.090 1704.770 ;
        RECT -22.670 1703.590 -21.490 1704.770 ;
        RECT -24.270 1701.990 -23.090 1703.170 ;
        RECT -22.670 1701.990 -21.490 1703.170 ;
        RECT -24.270 1523.590 -23.090 1524.770 ;
        RECT -22.670 1523.590 -21.490 1524.770 ;
        RECT -24.270 1521.990 -23.090 1523.170 ;
        RECT -22.670 1521.990 -21.490 1523.170 ;
        RECT -24.270 1343.590 -23.090 1344.770 ;
        RECT -22.670 1343.590 -21.490 1344.770 ;
        RECT -24.270 1341.990 -23.090 1343.170 ;
        RECT -22.670 1341.990 -21.490 1343.170 ;
        RECT -24.270 1163.590 -23.090 1164.770 ;
        RECT -22.670 1163.590 -21.490 1164.770 ;
        RECT -24.270 1161.990 -23.090 1163.170 ;
        RECT -22.670 1161.990 -21.490 1163.170 ;
        RECT -24.270 983.590 -23.090 984.770 ;
        RECT -22.670 983.590 -21.490 984.770 ;
        RECT -24.270 981.990 -23.090 983.170 ;
        RECT -22.670 981.990 -21.490 983.170 ;
        RECT -24.270 803.590 -23.090 804.770 ;
        RECT -22.670 803.590 -21.490 804.770 ;
        RECT -24.270 801.990 -23.090 803.170 ;
        RECT -22.670 801.990 -21.490 803.170 ;
        RECT -24.270 623.590 -23.090 624.770 ;
        RECT -22.670 623.590 -21.490 624.770 ;
        RECT -24.270 621.990 -23.090 623.170 ;
        RECT -22.670 621.990 -21.490 623.170 ;
        RECT -24.270 443.590 -23.090 444.770 ;
        RECT -22.670 443.590 -21.490 444.770 ;
        RECT -24.270 441.990 -23.090 443.170 ;
        RECT -22.670 441.990 -21.490 443.170 ;
        RECT -24.270 263.590 -23.090 264.770 ;
        RECT -22.670 263.590 -21.490 264.770 ;
        RECT -24.270 261.990 -23.090 263.170 ;
        RECT -22.670 261.990 -21.490 263.170 ;
        RECT -24.270 83.590 -23.090 84.770 ;
        RECT -22.670 83.590 -21.490 84.770 ;
        RECT -24.270 81.990 -23.090 83.170 ;
        RECT -22.670 81.990 -21.490 83.170 ;
        RECT -24.270 -17.310 -23.090 -16.130 ;
        RECT -22.670 -17.310 -21.490 -16.130 ;
        RECT -24.270 -18.910 -23.090 -17.730 ;
        RECT -22.670 -18.910 -21.490 -17.730 ;
        RECT 76.630 3537.410 77.810 3538.590 ;
        RECT 78.230 3537.410 79.410 3538.590 ;
        RECT 76.630 3535.810 77.810 3536.990 ;
        RECT 78.230 3535.810 79.410 3536.990 ;
        RECT 76.630 3503.590 77.810 3504.770 ;
        RECT 78.230 3503.590 79.410 3504.770 ;
        RECT 76.630 3501.990 77.810 3503.170 ;
        RECT 78.230 3501.990 79.410 3503.170 ;
        RECT 76.630 3323.590 77.810 3324.770 ;
        RECT 78.230 3323.590 79.410 3324.770 ;
        RECT 76.630 3321.990 77.810 3323.170 ;
        RECT 78.230 3321.990 79.410 3323.170 ;
        RECT 76.630 3143.590 77.810 3144.770 ;
        RECT 78.230 3143.590 79.410 3144.770 ;
        RECT 76.630 3141.990 77.810 3143.170 ;
        RECT 78.230 3141.990 79.410 3143.170 ;
        RECT 76.630 2963.590 77.810 2964.770 ;
        RECT 78.230 2963.590 79.410 2964.770 ;
        RECT 76.630 2961.990 77.810 2963.170 ;
        RECT 78.230 2961.990 79.410 2963.170 ;
        RECT 76.630 2783.590 77.810 2784.770 ;
        RECT 78.230 2783.590 79.410 2784.770 ;
        RECT 76.630 2781.990 77.810 2783.170 ;
        RECT 78.230 2781.990 79.410 2783.170 ;
        RECT 76.630 2603.590 77.810 2604.770 ;
        RECT 78.230 2603.590 79.410 2604.770 ;
        RECT 76.630 2601.990 77.810 2603.170 ;
        RECT 78.230 2601.990 79.410 2603.170 ;
        RECT 76.630 2423.590 77.810 2424.770 ;
        RECT 78.230 2423.590 79.410 2424.770 ;
        RECT 76.630 2421.990 77.810 2423.170 ;
        RECT 78.230 2421.990 79.410 2423.170 ;
        RECT 76.630 2243.590 77.810 2244.770 ;
        RECT 78.230 2243.590 79.410 2244.770 ;
        RECT 76.630 2241.990 77.810 2243.170 ;
        RECT 78.230 2241.990 79.410 2243.170 ;
        RECT 76.630 2063.590 77.810 2064.770 ;
        RECT 78.230 2063.590 79.410 2064.770 ;
        RECT 76.630 2061.990 77.810 2063.170 ;
        RECT 78.230 2061.990 79.410 2063.170 ;
        RECT 76.630 1883.590 77.810 1884.770 ;
        RECT 78.230 1883.590 79.410 1884.770 ;
        RECT 76.630 1881.990 77.810 1883.170 ;
        RECT 78.230 1881.990 79.410 1883.170 ;
        RECT 76.630 1703.590 77.810 1704.770 ;
        RECT 78.230 1703.590 79.410 1704.770 ;
        RECT 76.630 1701.990 77.810 1703.170 ;
        RECT 78.230 1701.990 79.410 1703.170 ;
        RECT 76.630 1523.590 77.810 1524.770 ;
        RECT 78.230 1523.590 79.410 1524.770 ;
        RECT 76.630 1521.990 77.810 1523.170 ;
        RECT 78.230 1521.990 79.410 1523.170 ;
        RECT 76.630 1343.590 77.810 1344.770 ;
        RECT 78.230 1343.590 79.410 1344.770 ;
        RECT 76.630 1341.990 77.810 1343.170 ;
        RECT 78.230 1341.990 79.410 1343.170 ;
        RECT 76.630 1163.590 77.810 1164.770 ;
        RECT 78.230 1163.590 79.410 1164.770 ;
        RECT 76.630 1161.990 77.810 1163.170 ;
        RECT 78.230 1161.990 79.410 1163.170 ;
        RECT 76.630 983.590 77.810 984.770 ;
        RECT 78.230 983.590 79.410 984.770 ;
        RECT 76.630 981.990 77.810 983.170 ;
        RECT 78.230 981.990 79.410 983.170 ;
        RECT 76.630 803.590 77.810 804.770 ;
        RECT 78.230 803.590 79.410 804.770 ;
        RECT 76.630 801.990 77.810 803.170 ;
        RECT 78.230 801.990 79.410 803.170 ;
        RECT 76.630 623.590 77.810 624.770 ;
        RECT 78.230 623.590 79.410 624.770 ;
        RECT 76.630 621.990 77.810 623.170 ;
        RECT 78.230 621.990 79.410 623.170 ;
        RECT 76.630 443.590 77.810 444.770 ;
        RECT 78.230 443.590 79.410 444.770 ;
        RECT 76.630 441.990 77.810 443.170 ;
        RECT 78.230 441.990 79.410 443.170 ;
        RECT 76.630 263.590 77.810 264.770 ;
        RECT 78.230 263.590 79.410 264.770 ;
        RECT 76.630 261.990 77.810 263.170 ;
        RECT 78.230 261.990 79.410 263.170 ;
        RECT 76.630 83.590 77.810 84.770 ;
        RECT 78.230 83.590 79.410 84.770 ;
        RECT 76.630 81.990 77.810 83.170 ;
        RECT 78.230 81.990 79.410 83.170 ;
        RECT 76.630 -17.310 77.810 -16.130 ;
        RECT 78.230 -17.310 79.410 -16.130 ;
        RECT 76.630 -18.910 77.810 -17.730 ;
        RECT 78.230 -18.910 79.410 -17.730 ;
        RECT 256.630 3537.410 257.810 3538.590 ;
        RECT 258.230 3537.410 259.410 3538.590 ;
        RECT 256.630 3535.810 257.810 3536.990 ;
        RECT 258.230 3535.810 259.410 3536.990 ;
        RECT 256.630 3503.590 257.810 3504.770 ;
        RECT 258.230 3503.590 259.410 3504.770 ;
        RECT 256.630 3501.990 257.810 3503.170 ;
        RECT 258.230 3501.990 259.410 3503.170 ;
        RECT 256.630 3323.590 257.810 3324.770 ;
        RECT 258.230 3323.590 259.410 3324.770 ;
        RECT 256.630 3321.990 257.810 3323.170 ;
        RECT 258.230 3321.990 259.410 3323.170 ;
        RECT 256.630 3143.590 257.810 3144.770 ;
        RECT 258.230 3143.590 259.410 3144.770 ;
        RECT 256.630 3141.990 257.810 3143.170 ;
        RECT 258.230 3141.990 259.410 3143.170 ;
        RECT 256.630 2963.590 257.810 2964.770 ;
        RECT 258.230 2963.590 259.410 2964.770 ;
        RECT 256.630 2961.990 257.810 2963.170 ;
        RECT 258.230 2961.990 259.410 2963.170 ;
        RECT 256.630 2783.590 257.810 2784.770 ;
        RECT 258.230 2783.590 259.410 2784.770 ;
        RECT 256.630 2781.990 257.810 2783.170 ;
        RECT 258.230 2781.990 259.410 2783.170 ;
        RECT 256.630 2603.590 257.810 2604.770 ;
        RECT 258.230 2603.590 259.410 2604.770 ;
        RECT 256.630 2601.990 257.810 2603.170 ;
        RECT 258.230 2601.990 259.410 2603.170 ;
        RECT 256.630 2423.590 257.810 2424.770 ;
        RECT 258.230 2423.590 259.410 2424.770 ;
        RECT 256.630 2421.990 257.810 2423.170 ;
        RECT 258.230 2421.990 259.410 2423.170 ;
        RECT 256.630 2243.590 257.810 2244.770 ;
        RECT 258.230 2243.590 259.410 2244.770 ;
        RECT 256.630 2241.990 257.810 2243.170 ;
        RECT 258.230 2241.990 259.410 2243.170 ;
        RECT 256.630 2063.590 257.810 2064.770 ;
        RECT 258.230 2063.590 259.410 2064.770 ;
        RECT 256.630 2061.990 257.810 2063.170 ;
        RECT 258.230 2061.990 259.410 2063.170 ;
        RECT 256.630 1883.590 257.810 1884.770 ;
        RECT 258.230 1883.590 259.410 1884.770 ;
        RECT 256.630 1881.990 257.810 1883.170 ;
        RECT 258.230 1881.990 259.410 1883.170 ;
        RECT 256.630 1703.590 257.810 1704.770 ;
        RECT 258.230 1703.590 259.410 1704.770 ;
        RECT 256.630 1701.990 257.810 1703.170 ;
        RECT 258.230 1701.990 259.410 1703.170 ;
        RECT 256.630 1523.590 257.810 1524.770 ;
        RECT 258.230 1523.590 259.410 1524.770 ;
        RECT 256.630 1521.990 257.810 1523.170 ;
        RECT 258.230 1521.990 259.410 1523.170 ;
        RECT 256.630 1343.590 257.810 1344.770 ;
        RECT 258.230 1343.590 259.410 1344.770 ;
        RECT 256.630 1341.990 257.810 1343.170 ;
        RECT 258.230 1341.990 259.410 1343.170 ;
        RECT 256.630 1163.590 257.810 1164.770 ;
        RECT 258.230 1163.590 259.410 1164.770 ;
        RECT 256.630 1161.990 257.810 1163.170 ;
        RECT 258.230 1161.990 259.410 1163.170 ;
        RECT 256.630 983.590 257.810 984.770 ;
        RECT 258.230 983.590 259.410 984.770 ;
        RECT 256.630 981.990 257.810 983.170 ;
        RECT 258.230 981.990 259.410 983.170 ;
        RECT 436.630 3537.410 437.810 3538.590 ;
        RECT 438.230 3537.410 439.410 3538.590 ;
        RECT 436.630 3535.810 437.810 3536.990 ;
        RECT 438.230 3535.810 439.410 3536.990 ;
        RECT 436.630 3503.590 437.810 3504.770 ;
        RECT 438.230 3503.590 439.410 3504.770 ;
        RECT 436.630 3501.990 437.810 3503.170 ;
        RECT 438.230 3501.990 439.410 3503.170 ;
        RECT 436.630 3323.590 437.810 3324.770 ;
        RECT 438.230 3323.590 439.410 3324.770 ;
        RECT 436.630 3321.990 437.810 3323.170 ;
        RECT 438.230 3321.990 439.410 3323.170 ;
        RECT 436.630 3143.590 437.810 3144.770 ;
        RECT 438.230 3143.590 439.410 3144.770 ;
        RECT 436.630 3141.990 437.810 3143.170 ;
        RECT 438.230 3141.990 439.410 3143.170 ;
        RECT 436.630 2963.590 437.810 2964.770 ;
        RECT 438.230 2963.590 439.410 2964.770 ;
        RECT 436.630 2961.990 437.810 2963.170 ;
        RECT 438.230 2961.990 439.410 2963.170 ;
        RECT 436.630 2783.590 437.810 2784.770 ;
        RECT 438.230 2783.590 439.410 2784.770 ;
        RECT 436.630 2781.990 437.810 2783.170 ;
        RECT 438.230 2781.990 439.410 2783.170 ;
        RECT 436.630 2603.590 437.810 2604.770 ;
        RECT 438.230 2603.590 439.410 2604.770 ;
        RECT 436.630 2601.990 437.810 2603.170 ;
        RECT 438.230 2601.990 439.410 2603.170 ;
        RECT 436.630 2423.590 437.810 2424.770 ;
        RECT 438.230 2423.590 439.410 2424.770 ;
        RECT 436.630 2421.990 437.810 2423.170 ;
        RECT 438.230 2421.990 439.410 2423.170 ;
        RECT 436.630 2243.590 437.810 2244.770 ;
        RECT 438.230 2243.590 439.410 2244.770 ;
        RECT 436.630 2241.990 437.810 2243.170 ;
        RECT 438.230 2241.990 439.410 2243.170 ;
        RECT 436.630 2063.590 437.810 2064.770 ;
        RECT 438.230 2063.590 439.410 2064.770 ;
        RECT 436.630 2061.990 437.810 2063.170 ;
        RECT 438.230 2061.990 439.410 2063.170 ;
        RECT 436.630 1883.590 437.810 1884.770 ;
        RECT 438.230 1883.590 439.410 1884.770 ;
        RECT 436.630 1881.990 437.810 1883.170 ;
        RECT 438.230 1881.990 439.410 1883.170 ;
        RECT 436.630 1703.590 437.810 1704.770 ;
        RECT 438.230 1703.590 439.410 1704.770 ;
        RECT 436.630 1701.990 437.810 1703.170 ;
        RECT 438.230 1701.990 439.410 1703.170 ;
        RECT 436.630 1523.590 437.810 1524.770 ;
        RECT 438.230 1523.590 439.410 1524.770 ;
        RECT 436.630 1521.990 437.810 1523.170 ;
        RECT 438.230 1521.990 439.410 1523.170 ;
        RECT 436.630 1343.590 437.810 1344.770 ;
        RECT 438.230 1343.590 439.410 1344.770 ;
        RECT 436.630 1341.990 437.810 1343.170 ;
        RECT 438.230 1341.990 439.410 1343.170 ;
        RECT 436.630 1163.590 437.810 1164.770 ;
        RECT 438.230 1163.590 439.410 1164.770 ;
        RECT 436.630 1161.990 437.810 1163.170 ;
        RECT 438.230 1161.990 439.410 1163.170 ;
        RECT 436.630 983.590 437.810 984.770 ;
        RECT 438.230 983.590 439.410 984.770 ;
        RECT 436.630 981.990 437.810 983.170 ;
        RECT 438.230 981.990 439.410 983.170 ;
        RECT 616.630 3537.410 617.810 3538.590 ;
        RECT 618.230 3537.410 619.410 3538.590 ;
        RECT 616.630 3535.810 617.810 3536.990 ;
        RECT 618.230 3535.810 619.410 3536.990 ;
        RECT 616.630 3503.590 617.810 3504.770 ;
        RECT 618.230 3503.590 619.410 3504.770 ;
        RECT 616.630 3501.990 617.810 3503.170 ;
        RECT 618.230 3501.990 619.410 3503.170 ;
        RECT 616.630 3323.590 617.810 3324.770 ;
        RECT 618.230 3323.590 619.410 3324.770 ;
        RECT 616.630 3321.990 617.810 3323.170 ;
        RECT 618.230 3321.990 619.410 3323.170 ;
        RECT 616.630 3143.590 617.810 3144.770 ;
        RECT 618.230 3143.590 619.410 3144.770 ;
        RECT 616.630 3141.990 617.810 3143.170 ;
        RECT 618.230 3141.990 619.410 3143.170 ;
        RECT 616.630 2963.590 617.810 2964.770 ;
        RECT 618.230 2963.590 619.410 2964.770 ;
        RECT 616.630 2961.990 617.810 2963.170 ;
        RECT 618.230 2961.990 619.410 2963.170 ;
        RECT 616.630 2783.590 617.810 2784.770 ;
        RECT 618.230 2783.590 619.410 2784.770 ;
        RECT 616.630 2781.990 617.810 2783.170 ;
        RECT 618.230 2781.990 619.410 2783.170 ;
        RECT 616.630 2603.590 617.810 2604.770 ;
        RECT 618.230 2603.590 619.410 2604.770 ;
        RECT 616.630 2601.990 617.810 2603.170 ;
        RECT 618.230 2601.990 619.410 2603.170 ;
        RECT 616.630 2423.590 617.810 2424.770 ;
        RECT 618.230 2423.590 619.410 2424.770 ;
        RECT 616.630 2421.990 617.810 2423.170 ;
        RECT 618.230 2421.990 619.410 2423.170 ;
        RECT 616.630 2243.590 617.810 2244.770 ;
        RECT 618.230 2243.590 619.410 2244.770 ;
        RECT 616.630 2241.990 617.810 2243.170 ;
        RECT 618.230 2241.990 619.410 2243.170 ;
        RECT 616.630 2063.590 617.810 2064.770 ;
        RECT 618.230 2063.590 619.410 2064.770 ;
        RECT 616.630 2061.990 617.810 2063.170 ;
        RECT 618.230 2061.990 619.410 2063.170 ;
        RECT 616.630 1883.590 617.810 1884.770 ;
        RECT 618.230 1883.590 619.410 1884.770 ;
        RECT 616.630 1881.990 617.810 1883.170 ;
        RECT 618.230 1881.990 619.410 1883.170 ;
        RECT 616.630 1703.590 617.810 1704.770 ;
        RECT 618.230 1703.590 619.410 1704.770 ;
        RECT 616.630 1701.990 617.810 1703.170 ;
        RECT 618.230 1701.990 619.410 1703.170 ;
        RECT 616.630 1523.590 617.810 1524.770 ;
        RECT 618.230 1523.590 619.410 1524.770 ;
        RECT 616.630 1521.990 617.810 1523.170 ;
        RECT 618.230 1521.990 619.410 1523.170 ;
        RECT 616.630 1343.590 617.810 1344.770 ;
        RECT 618.230 1343.590 619.410 1344.770 ;
        RECT 616.630 1341.990 617.810 1343.170 ;
        RECT 618.230 1341.990 619.410 1343.170 ;
        RECT 616.630 1163.590 617.810 1164.770 ;
        RECT 618.230 1163.590 619.410 1164.770 ;
        RECT 616.630 1161.990 617.810 1163.170 ;
        RECT 618.230 1161.990 619.410 1163.170 ;
        RECT 616.630 983.590 617.810 984.770 ;
        RECT 618.230 983.590 619.410 984.770 ;
        RECT 616.630 981.990 617.810 983.170 ;
        RECT 618.230 981.990 619.410 983.170 ;
        RECT 796.630 3537.410 797.810 3538.590 ;
        RECT 798.230 3537.410 799.410 3538.590 ;
        RECT 796.630 3535.810 797.810 3536.990 ;
        RECT 798.230 3535.810 799.410 3536.990 ;
        RECT 796.630 3503.590 797.810 3504.770 ;
        RECT 798.230 3503.590 799.410 3504.770 ;
        RECT 796.630 3501.990 797.810 3503.170 ;
        RECT 798.230 3501.990 799.410 3503.170 ;
        RECT 796.630 3323.590 797.810 3324.770 ;
        RECT 798.230 3323.590 799.410 3324.770 ;
        RECT 796.630 3321.990 797.810 3323.170 ;
        RECT 798.230 3321.990 799.410 3323.170 ;
        RECT 796.630 3143.590 797.810 3144.770 ;
        RECT 798.230 3143.590 799.410 3144.770 ;
        RECT 796.630 3141.990 797.810 3143.170 ;
        RECT 798.230 3141.990 799.410 3143.170 ;
        RECT 796.630 2963.590 797.810 2964.770 ;
        RECT 798.230 2963.590 799.410 2964.770 ;
        RECT 796.630 2961.990 797.810 2963.170 ;
        RECT 798.230 2961.990 799.410 2963.170 ;
        RECT 796.630 2783.590 797.810 2784.770 ;
        RECT 798.230 2783.590 799.410 2784.770 ;
        RECT 796.630 2781.990 797.810 2783.170 ;
        RECT 798.230 2781.990 799.410 2783.170 ;
        RECT 796.630 2603.590 797.810 2604.770 ;
        RECT 798.230 2603.590 799.410 2604.770 ;
        RECT 796.630 2601.990 797.810 2603.170 ;
        RECT 798.230 2601.990 799.410 2603.170 ;
        RECT 796.630 2423.590 797.810 2424.770 ;
        RECT 798.230 2423.590 799.410 2424.770 ;
        RECT 796.630 2421.990 797.810 2423.170 ;
        RECT 798.230 2421.990 799.410 2423.170 ;
        RECT 796.630 2243.590 797.810 2244.770 ;
        RECT 798.230 2243.590 799.410 2244.770 ;
        RECT 796.630 2241.990 797.810 2243.170 ;
        RECT 798.230 2241.990 799.410 2243.170 ;
        RECT 796.630 2063.590 797.810 2064.770 ;
        RECT 798.230 2063.590 799.410 2064.770 ;
        RECT 796.630 2061.990 797.810 2063.170 ;
        RECT 798.230 2061.990 799.410 2063.170 ;
        RECT 796.630 1883.590 797.810 1884.770 ;
        RECT 798.230 1883.590 799.410 1884.770 ;
        RECT 796.630 1881.990 797.810 1883.170 ;
        RECT 798.230 1881.990 799.410 1883.170 ;
        RECT 796.630 1703.590 797.810 1704.770 ;
        RECT 798.230 1703.590 799.410 1704.770 ;
        RECT 796.630 1701.990 797.810 1703.170 ;
        RECT 798.230 1701.990 799.410 1703.170 ;
        RECT 796.630 1523.590 797.810 1524.770 ;
        RECT 798.230 1523.590 799.410 1524.770 ;
        RECT 796.630 1521.990 797.810 1523.170 ;
        RECT 798.230 1521.990 799.410 1523.170 ;
        RECT 796.630 1343.590 797.810 1344.770 ;
        RECT 798.230 1343.590 799.410 1344.770 ;
        RECT 796.630 1341.990 797.810 1343.170 ;
        RECT 798.230 1341.990 799.410 1343.170 ;
        RECT 796.630 1163.590 797.810 1164.770 ;
        RECT 798.230 1163.590 799.410 1164.770 ;
        RECT 796.630 1161.990 797.810 1163.170 ;
        RECT 798.230 1161.990 799.410 1163.170 ;
        RECT 796.630 983.590 797.810 984.770 ;
        RECT 798.230 983.590 799.410 984.770 ;
        RECT 796.630 981.990 797.810 983.170 ;
        RECT 798.230 981.990 799.410 983.170 ;
        RECT 256.630 803.590 257.810 804.770 ;
        RECT 258.230 803.590 259.410 804.770 ;
        RECT 256.630 801.990 257.810 803.170 ;
        RECT 258.230 801.990 259.410 803.170 ;
        RECT 256.630 623.590 257.810 624.770 ;
        RECT 258.230 623.590 259.410 624.770 ;
        RECT 256.630 621.990 257.810 623.170 ;
        RECT 258.230 621.990 259.410 623.170 ;
        RECT 796.630 803.590 797.810 804.770 ;
        RECT 798.230 803.590 799.410 804.770 ;
        RECT 796.630 801.990 797.810 803.170 ;
        RECT 798.230 801.990 799.410 803.170 ;
        RECT 796.630 623.590 797.810 624.770 ;
        RECT 798.230 623.590 799.410 624.770 ;
        RECT 796.630 621.990 797.810 623.170 ;
        RECT 798.230 621.990 799.410 623.170 ;
        RECT 256.630 443.590 257.810 444.770 ;
        RECT 258.230 443.590 259.410 444.770 ;
        RECT 256.630 441.990 257.810 443.170 ;
        RECT 258.230 441.990 259.410 443.170 ;
        RECT 256.630 263.590 257.810 264.770 ;
        RECT 258.230 263.590 259.410 264.770 ;
        RECT 256.630 261.990 257.810 263.170 ;
        RECT 258.230 261.990 259.410 263.170 ;
        RECT 256.630 83.590 257.810 84.770 ;
        RECT 258.230 83.590 259.410 84.770 ;
        RECT 256.630 81.990 257.810 83.170 ;
        RECT 258.230 81.990 259.410 83.170 ;
        RECT 256.630 -17.310 257.810 -16.130 ;
        RECT 258.230 -17.310 259.410 -16.130 ;
        RECT 256.630 -18.910 257.810 -17.730 ;
        RECT 258.230 -18.910 259.410 -17.730 ;
        RECT 436.630 443.590 437.810 444.770 ;
        RECT 438.230 443.590 439.410 444.770 ;
        RECT 436.630 441.990 437.810 443.170 ;
        RECT 438.230 441.990 439.410 443.170 ;
        RECT 436.630 263.590 437.810 264.770 ;
        RECT 438.230 263.590 439.410 264.770 ;
        RECT 436.630 261.990 437.810 263.170 ;
        RECT 438.230 261.990 439.410 263.170 ;
        RECT 436.630 83.590 437.810 84.770 ;
        RECT 438.230 83.590 439.410 84.770 ;
        RECT 436.630 81.990 437.810 83.170 ;
        RECT 438.230 81.990 439.410 83.170 ;
        RECT 436.630 -17.310 437.810 -16.130 ;
        RECT 438.230 -17.310 439.410 -16.130 ;
        RECT 436.630 -18.910 437.810 -17.730 ;
        RECT 438.230 -18.910 439.410 -17.730 ;
        RECT 616.630 443.590 617.810 444.770 ;
        RECT 618.230 443.590 619.410 444.770 ;
        RECT 616.630 441.990 617.810 443.170 ;
        RECT 618.230 441.990 619.410 443.170 ;
        RECT 616.630 263.590 617.810 264.770 ;
        RECT 618.230 263.590 619.410 264.770 ;
        RECT 616.630 261.990 617.810 263.170 ;
        RECT 618.230 261.990 619.410 263.170 ;
        RECT 616.630 83.590 617.810 84.770 ;
        RECT 618.230 83.590 619.410 84.770 ;
        RECT 616.630 81.990 617.810 83.170 ;
        RECT 618.230 81.990 619.410 83.170 ;
        RECT 616.630 -17.310 617.810 -16.130 ;
        RECT 618.230 -17.310 619.410 -16.130 ;
        RECT 616.630 -18.910 617.810 -17.730 ;
        RECT 618.230 -18.910 619.410 -17.730 ;
        RECT 796.630 443.590 797.810 444.770 ;
        RECT 798.230 443.590 799.410 444.770 ;
        RECT 796.630 441.990 797.810 443.170 ;
        RECT 798.230 441.990 799.410 443.170 ;
        RECT 796.630 263.590 797.810 264.770 ;
        RECT 798.230 263.590 799.410 264.770 ;
        RECT 796.630 261.990 797.810 263.170 ;
        RECT 798.230 261.990 799.410 263.170 ;
        RECT 796.630 83.590 797.810 84.770 ;
        RECT 798.230 83.590 799.410 84.770 ;
        RECT 796.630 81.990 797.810 83.170 ;
        RECT 798.230 81.990 799.410 83.170 ;
        RECT 796.630 -17.310 797.810 -16.130 ;
        RECT 798.230 -17.310 799.410 -16.130 ;
        RECT 796.630 -18.910 797.810 -17.730 ;
        RECT 798.230 -18.910 799.410 -17.730 ;
        RECT 976.630 3537.410 977.810 3538.590 ;
        RECT 978.230 3537.410 979.410 3538.590 ;
        RECT 976.630 3535.810 977.810 3536.990 ;
        RECT 978.230 3535.810 979.410 3536.990 ;
        RECT 976.630 3503.590 977.810 3504.770 ;
        RECT 978.230 3503.590 979.410 3504.770 ;
        RECT 976.630 3501.990 977.810 3503.170 ;
        RECT 978.230 3501.990 979.410 3503.170 ;
        RECT 976.630 3323.590 977.810 3324.770 ;
        RECT 978.230 3323.590 979.410 3324.770 ;
        RECT 976.630 3321.990 977.810 3323.170 ;
        RECT 978.230 3321.990 979.410 3323.170 ;
        RECT 976.630 3143.590 977.810 3144.770 ;
        RECT 978.230 3143.590 979.410 3144.770 ;
        RECT 976.630 3141.990 977.810 3143.170 ;
        RECT 978.230 3141.990 979.410 3143.170 ;
        RECT 976.630 2963.590 977.810 2964.770 ;
        RECT 978.230 2963.590 979.410 2964.770 ;
        RECT 976.630 2961.990 977.810 2963.170 ;
        RECT 978.230 2961.990 979.410 2963.170 ;
        RECT 976.630 2783.590 977.810 2784.770 ;
        RECT 978.230 2783.590 979.410 2784.770 ;
        RECT 976.630 2781.990 977.810 2783.170 ;
        RECT 978.230 2781.990 979.410 2783.170 ;
        RECT 976.630 2603.590 977.810 2604.770 ;
        RECT 978.230 2603.590 979.410 2604.770 ;
        RECT 976.630 2601.990 977.810 2603.170 ;
        RECT 978.230 2601.990 979.410 2603.170 ;
        RECT 976.630 2423.590 977.810 2424.770 ;
        RECT 978.230 2423.590 979.410 2424.770 ;
        RECT 976.630 2421.990 977.810 2423.170 ;
        RECT 978.230 2421.990 979.410 2423.170 ;
        RECT 976.630 2243.590 977.810 2244.770 ;
        RECT 978.230 2243.590 979.410 2244.770 ;
        RECT 976.630 2241.990 977.810 2243.170 ;
        RECT 978.230 2241.990 979.410 2243.170 ;
        RECT 976.630 2063.590 977.810 2064.770 ;
        RECT 978.230 2063.590 979.410 2064.770 ;
        RECT 976.630 2061.990 977.810 2063.170 ;
        RECT 978.230 2061.990 979.410 2063.170 ;
        RECT 976.630 1883.590 977.810 1884.770 ;
        RECT 978.230 1883.590 979.410 1884.770 ;
        RECT 976.630 1881.990 977.810 1883.170 ;
        RECT 978.230 1881.990 979.410 1883.170 ;
        RECT 976.630 1703.590 977.810 1704.770 ;
        RECT 978.230 1703.590 979.410 1704.770 ;
        RECT 976.630 1701.990 977.810 1703.170 ;
        RECT 978.230 1701.990 979.410 1703.170 ;
        RECT 976.630 1523.590 977.810 1524.770 ;
        RECT 978.230 1523.590 979.410 1524.770 ;
        RECT 976.630 1521.990 977.810 1523.170 ;
        RECT 978.230 1521.990 979.410 1523.170 ;
        RECT 976.630 1343.590 977.810 1344.770 ;
        RECT 978.230 1343.590 979.410 1344.770 ;
        RECT 976.630 1341.990 977.810 1343.170 ;
        RECT 978.230 1341.990 979.410 1343.170 ;
        RECT 976.630 1163.590 977.810 1164.770 ;
        RECT 978.230 1163.590 979.410 1164.770 ;
        RECT 976.630 1161.990 977.810 1163.170 ;
        RECT 978.230 1161.990 979.410 1163.170 ;
        RECT 976.630 983.590 977.810 984.770 ;
        RECT 978.230 983.590 979.410 984.770 ;
        RECT 976.630 981.990 977.810 983.170 ;
        RECT 978.230 981.990 979.410 983.170 ;
        RECT 976.630 803.590 977.810 804.770 ;
        RECT 978.230 803.590 979.410 804.770 ;
        RECT 976.630 801.990 977.810 803.170 ;
        RECT 978.230 801.990 979.410 803.170 ;
        RECT 976.630 623.590 977.810 624.770 ;
        RECT 978.230 623.590 979.410 624.770 ;
        RECT 976.630 621.990 977.810 623.170 ;
        RECT 978.230 621.990 979.410 623.170 ;
        RECT 976.630 443.590 977.810 444.770 ;
        RECT 978.230 443.590 979.410 444.770 ;
        RECT 976.630 441.990 977.810 443.170 ;
        RECT 978.230 441.990 979.410 443.170 ;
        RECT 976.630 263.590 977.810 264.770 ;
        RECT 978.230 263.590 979.410 264.770 ;
        RECT 976.630 261.990 977.810 263.170 ;
        RECT 978.230 261.990 979.410 263.170 ;
        RECT 976.630 83.590 977.810 84.770 ;
        RECT 978.230 83.590 979.410 84.770 ;
        RECT 976.630 81.990 977.810 83.170 ;
        RECT 978.230 81.990 979.410 83.170 ;
        RECT 976.630 -17.310 977.810 -16.130 ;
        RECT 978.230 -17.310 979.410 -16.130 ;
        RECT 976.630 -18.910 977.810 -17.730 ;
        RECT 978.230 -18.910 979.410 -17.730 ;
        RECT 1156.630 3537.410 1157.810 3538.590 ;
        RECT 1158.230 3537.410 1159.410 3538.590 ;
        RECT 1156.630 3535.810 1157.810 3536.990 ;
        RECT 1158.230 3535.810 1159.410 3536.990 ;
        RECT 1156.630 3503.590 1157.810 3504.770 ;
        RECT 1158.230 3503.590 1159.410 3504.770 ;
        RECT 1156.630 3501.990 1157.810 3503.170 ;
        RECT 1158.230 3501.990 1159.410 3503.170 ;
        RECT 1156.630 3323.590 1157.810 3324.770 ;
        RECT 1158.230 3323.590 1159.410 3324.770 ;
        RECT 1156.630 3321.990 1157.810 3323.170 ;
        RECT 1158.230 3321.990 1159.410 3323.170 ;
        RECT 1156.630 3143.590 1157.810 3144.770 ;
        RECT 1158.230 3143.590 1159.410 3144.770 ;
        RECT 1156.630 3141.990 1157.810 3143.170 ;
        RECT 1158.230 3141.990 1159.410 3143.170 ;
        RECT 1156.630 2963.590 1157.810 2964.770 ;
        RECT 1158.230 2963.590 1159.410 2964.770 ;
        RECT 1156.630 2961.990 1157.810 2963.170 ;
        RECT 1158.230 2961.990 1159.410 2963.170 ;
        RECT 1156.630 2783.590 1157.810 2784.770 ;
        RECT 1158.230 2783.590 1159.410 2784.770 ;
        RECT 1156.630 2781.990 1157.810 2783.170 ;
        RECT 1158.230 2781.990 1159.410 2783.170 ;
        RECT 1156.630 2603.590 1157.810 2604.770 ;
        RECT 1158.230 2603.590 1159.410 2604.770 ;
        RECT 1156.630 2601.990 1157.810 2603.170 ;
        RECT 1158.230 2601.990 1159.410 2603.170 ;
        RECT 1156.630 2423.590 1157.810 2424.770 ;
        RECT 1158.230 2423.590 1159.410 2424.770 ;
        RECT 1156.630 2421.990 1157.810 2423.170 ;
        RECT 1158.230 2421.990 1159.410 2423.170 ;
        RECT 1156.630 2243.590 1157.810 2244.770 ;
        RECT 1158.230 2243.590 1159.410 2244.770 ;
        RECT 1156.630 2241.990 1157.810 2243.170 ;
        RECT 1158.230 2241.990 1159.410 2243.170 ;
        RECT 1156.630 2063.590 1157.810 2064.770 ;
        RECT 1158.230 2063.590 1159.410 2064.770 ;
        RECT 1156.630 2061.990 1157.810 2063.170 ;
        RECT 1158.230 2061.990 1159.410 2063.170 ;
        RECT 1156.630 1883.590 1157.810 1884.770 ;
        RECT 1158.230 1883.590 1159.410 1884.770 ;
        RECT 1156.630 1881.990 1157.810 1883.170 ;
        RECT 1158.230 1881.990 1159.410 1883.170 ;
        RECT 1156.630 1703.590 1157.810 1704.770 ;
        RECT 1158.230 1703.590 1159.410 1704.770 ;
        RECT 1156.630 1701.990 1157.810 1703.170 ;
        RECT 1158.230 1701.990 1159.410 1703.170 ;
        RECT 1156.630 1523.590 1157.810 1524.770 ;
        RECT 1158.230 1523.590 1159.410 1524.770 ;
        RECT 1156.630 1521.990 1157.810 1523.170 ;
        RECT 1158.230 1521.990 1159.410 1523.170 ;
        RECT 1156.630 1343.590 1157.810 1344.770 ;
        RECT 1158.230 1343.590 1159.410 1344.770 ;
        RECT 1156.630 1341.990 1157.810 1343.170 ;
        RECT 1158.230 1341.990 1159.410 1343.170 ;
        RECT 1156.630 1163.590 1157.810 1164.770 ;
        RECT 1158.230 1163.590 1159.410 1164.770 ;
        RECT 1156.630 1161.990 1157.810 1163.170 ;
        RECT 1158.230 1161.990 1159.410 1163.170 ;
        RECT 1156.630 983.590 1157.810 984.770 ;
        RECT 1158.230 983.590 1159.410 984.770 ;
        RECT 1156.630 981.990 1157.810 983.170 ;
        RECT 1158.230 981.990 1159.410 983.170 ;
        RECT 1156.630 803.590 1157.810 804.770 ;
        RECT 1158.230 803.590 1159.410 804.770 ;
        RECT 1156.630 801.990 1157.810 803.170 ;
        RECT 1158.230 801.990 1159.410 803.170 ;
        RECT 1156.630 623.590 1157.810 624.770 ;
        RECT 1158.230 623.590 1159.410 624.770 ;
        RECT 1156.630 621.990 1157.810 623.170 ;
        RECT 1158.230 621.990 1159.410 623.170 ;
        RECT 1156.630 443.590 1157.810 444.770 ;
        RECT 1158.230 443.590 1159.410 444.770 ;
        RECT 1156.630 441.990 1157.810 443.170 ;
        RECT 1158.230 441.990 1159.410 443.170 ;
        RECT 1156.630 263.590 1157.810 264.770 ;
        RECT 1158.230 263.590 1159.410 264.770 ;
        RECT 1156.630 261.990 1157.810 263.170 ;
        RECT 1158.230 261.990 1159.410 263.170 ;
        RECT 1156.630 83.590 1157.810 84.770 ;
        RECT 1158.230 83.590 1159.410 84.770 ;
        RECT 1156.630 81.990 1157.810 83.170 ;
        RECT 1158.230 81.990 1159.410 83.170 ;
        RECT 1156.630 -17.310 1157.810 -16.130 ;
        RECT 1158.230 -17.310 1159.410 -16.130 ;
        RECT 1156.630 -18.910 1157.810 -17.730 ;
        RECT 1158.230 -18.910 1159.410 -17.730 ;
        RECT 1336.630 3537.410 1337.810 3538.590 ;
        RECT 1338.230 3537.410 1339.410 3538.590 ;
        RECT 1336.630 3535.810 1337.810 3536.990 ;
        RECT 1338.230 3535.810 1339.410 3536.990 ;
        RECT 1336.630 3503.590 1337.810 3504.770 ;
        RECT 1338.230 3503.590 1339.410 3504.770 ;
        RECT 1336.630 3501.990 1337.810 3503.170 ;
        RECT 1338.230 3501.990 1339.410 3503.170 ;
        RECT 1336.630 3323.590 1337.810 3324.770 ;
        RECT 1338.230 3323.590 1339.410 3324.770 ;
        RECT 1336.630 3321.990 1337.810 3323.170 ;
        RECT 1338.230 3321.990 1339.410 3323.170 ;
        RECT 1336.630 3143.590 1337.810 3144.770 ;
        RECT 1338.230 3143.590 1339.410 3144.770 ;
        RECT 1336.630 3141.990 1337.810 3143.170 ;
        RECT 1338.230 3141.990 1339.410 3143.170 ;
        RECT 1336.630 2963.590 1337.810 2964.770 ;
        RECT 1338.230 2963.590 1339.410 2964.770 ;
        RECT 1336.630 2961.990 1337.810 2963.170 ;
        RECT 1338.230 2961.990 1339.410 2963.170 ;
        RECT 1336.630 2783.590 1337.810 2784.770 ;
        RECT 1338.230 2783.590 1339.410 2784.770 ;
        RECT 1336.630 2781.990 1337.810 2783.170 ;
        RECT 1338.230 2781.990 1339.410 2783.170 ;
        RECT 1336.630 2603.590 1337.810 2604.770 ;
        RECT 1338.230 2603.590 1339.410 2604.770 ;
        RECT 1336.630 2601.990 1337.810 2603.170 ;
        RECT 1338.230 2601.990 1339.410 2603.170 ;
        RECT 1336.630 2423.590 1337.810 2424.770 ;
        RECT 1338.230 2423.590 1339.410 2424.770 ;
        RECT 1336.630 2421.990 1337.810 2423.170 ;
        RECT 1338.230 2421.990 1339.410 2423.170 ;
        RECT 1336.630 2243.590 1337.810 2244.770 ;
        RECT 1338.230 2243.590 1339.410 2244.770 ;
        RECT 1336.630 2241.990 1337.810 2243.170 ;
        RECT 1338.230 2241.990 1339.410 2243.170 ;
        RECT 1336.630 2063.590 1337.810 2064.770 ;
        RECT 1338.230 2063.590 1339.410 2064.770 ;
        RECT 1336.630 2061.990 1337.810 2063.170 ;
        RECT 1338.230 2061.990 1339.410 2063.170 ;
        RECT 1336.630 1883.590 1337.810 1884.770 ;
        RECT 1338.230 1883.590 1339.410 1884.770 ;
        RECT 1336.630 1881.990 1337.810 1883.170 ;
        RECT 1338.230 1881.990 1339.410 1883.170 ;
        RECT 1336.630 1703.590 1337.810 1704.770 ;
        RECT 1338.230 1703.590 1339.410 1704.770 ;
        RECT 1336.630 1701.990 1337.810 1703.170 ;
        RECT 1338.230 1701.990 1339.410 1703.170 ;
        RECT 1336.630 1523.590 1337.810 1524.770 ;
        RECT 1338.230 1523.590 1339.410 1524.770 ;
        RECT 1336.630 1521.990 1337.810 1523.170 ;
        RECT 1338.230 1521.990 1339.410 1523.170 ;
        RECT 1336.630 1343.590 1337.810 1344.770 ;
        RECT 1338.230 1343.590 1339.410 1344.770 ;
        RECT 1336.630 1341.990 1337.810 1343.170 ;
        RECT 1338.230 1341.990 1339.410 1343.170 ;
        RECT 1336.630 1163.590 1337.810 1164.770 ;
        RECT 1338.230 1163.590 1339.410 1164.770 ;
        RECT 1336.630 1161.990 1337.810 1163.170 ;
        RECT 1338.230 1161.990 1339.410 1163.170 ;
        RECT 1336.630 983.590 1337.810 984.770 ;
        RECT 1338.230 983.590 1339.410 984.770 ;
        RECT 1336.630 981.990 1337.810 983.170 ;
        RECT 1338.230 981.990 1339.410 983.170 ;
        RECT 1336.630 803.590 1337.810 804.770 ;
        RECT 1338.230 803.590 1339.410 804.770 ;
        RECT 1336.630 801.990 1337.810 803.170 ;
        RECT 1338.230 801.990 1339.410 803.170 ;
        RECT 1336.630 623.590 1337.810 624.770 ;
        RECT 1338.230 623.590 1339.410 624.770 ;
        RECT 1336.630 621.990 1337.810 623.170 ;
        RECT 1338.230 621.990 1339.410 623.170 ;
        RECT 1336.630 443.590 1337.810 444.770 ;
        RECT 1338.230 443.590 1339.410 444.770 ;
        RECT 1336.630 441.990 1337.810 443.170 ;
        RECT 1338.230 441.990 1339.410 443.170 ;
        RECT 1336.630 263.590 1337.810 264.770 ;
        RECT 1338.230 263.590 1339.410 264.770 ;
        RECT 1336.630 261.990 1337.810 263.170 ;
        RECT 1338.230 261.990 1339.410 263.170 ;
        RECT 1336.630 83.590 1337.810 84.770 ;
        RECT 1338.230 83.590 1339.410 84.770 ;
        RECT 1336.630 81.990 1337.810 83.170 ;
        RECT 1338.230 81.990 1339.410 83.170 ;
        RECT 1336.630 -17.310 1337.810 -16.130 ;
        RECT 1338.230 -17.310 1339.410 -16.130 ;
        RECT 1336.630 -18.910 1337.810 -17.730 ;
        RECT 1338.230 -18.910 1339.410 -17.730 ;
        RECT 1516.630 3537.410 1517.810 3538.590 ;
        RECT 1518.230 3537.410 1519.410 3538.590 ;
        RECT 1516.630 3535.810 1517.810 3536.990 ;
        RECT 1518.230 3535.810 1519.410 3536.990 ;
        RECT 1516.630 3503.590 1517.810 3504.770 ;
        RECT 1518.230 3503.590 1519.410 3504.770 ;
        RECT 1516.630 3501.990 1517.810 3503.170 ;
        RECT 1518.230 3501.990 1519.410 3503.170 ;
        RECT 1516.630 3323.590 1517.810 3324.770 ;
        RECT 1518.230 3323.590 1519.410 3324.770 ;
        RECT 1516.630 3321.990 1517.810 3323.170 ;
        RECT 1518.230 3321.990 1519.410 3323.170 ;
        RECT 1516.630 3143.590 1517.810 3144.770 ;
        RECT 1518.230 3143.590 1519.410 3144.770 ;
        RECT 1516.630 3141.990 1517.810 3143.170 ;
        RECT 1518.230 3141.990 1519.410 3143.170 ;
        RECT 1516.630 2963.590 1517.810 2964.770 ;
        RECT 1518.230 2963.590 1519.410 2964.770 ;
        RECT 1516.630 2961.990 1517.810 2963.170 ;
        RECT 1518.230 2961.990 1519.410 2963.170 ;
        RECT 1516.630 2783.590 1517.810 2784.770 ;
        RECT 1518.230 2783.590 1519.410 2784.770 ;
        RECT 1516.630 2781.990 1517.810 2783.170 ;
        RECT 1518.230 2781.990 1519.410 2783.170 ;
        RECT 1516.630 2603.590 1517.810 2604.770 ;
        RECT 1518.230 2603.590 1519.410 2604.770 ;
        RECT 1516.630 2601.990 1517.810 2603.170 ;
        RECT 1518.230 2601.990 1519.410 2603.170 ;
        RECT 1516.630 2423.590 1517.810 2424.770 ;
        RECT 1518.230 2423.590 1519.410 2424.770 ;
        RECT 1516.630 2421.990 1517.810 2423.170 ;
        RECT 1518.230 2421.990 1519.410 2423.170 ;
        RECT 1516.630 2243.590 1517.810 2244.770 ;
        RECT 1518.230 2243.590 1519.410 2244.770 ;
        RECT 1516.630 2241.990 1517.810 2243.170 ;
        RECT 1518.230 2241.990 1519.410 2243.170 ;
        RECT 1516.630 2063.590 1517.810 2064.770 ;
        RECT 1518.230 2063.590 1519.410 2064.770 ;
        RECT 1516.630 2061.990 1517.810 2063.170 ;
        RECT 1518.230 2061.990 1519.410 2063.170 ;
        RECT 1516.630 1883.590 1517.810 1884.770 ;
        RECT 1518.230 1883.590 1519.410 1884.770 ;
        RECT 1516.630 1881.990 1517.810 1883.170 ;
        RECT 1518.230 1881.990 1519.410 1883.170 ;
        RECT 1516.630 1703.590 1517.810 1704.770 ;
        RECT 1518.230 1703.590 1519.410 1704.770 ;
        RECT 1516.630 1701.990 1517.810 1703.170 ;
        RECT 1518.230 1701.990 1519.410 1703.170 ;
        RECT 1516.630 1523.590 1517.810 1524.770 ;
        RECT 1518.230 1523.590 1519.410 1524.770 ;
        RECT 1516.630 1521.990 1517.810 1523.170 ;
        RECT 1518.230 1521.990 1519.410 1523.170 ;
        RECT 1516.630 1343.590 1517.810 1344.770 ;
        RECT 1518.230 1343.590 1519.410 1344.770 ;
        RECT 1516.630 1341.990 1517.810 1343.170 ;
        RECT 1518.230 1341.990 1519.410 1343.170 ;
        RECT 1516.630 1163.590 1517.810 1164.770 ;
        RECT 1518.230 1163.590 1519.410 1164.770 ;
        RECT 1516.630 1161.990 1517.810 1163.170 ;
        RECT 1518.230 1161.990 1519.410 1163.170 ;
        RECT 1516.630 983.590 1517.810 984.770 ;
        RECT 1518.230 983.590 1519.410 984.770 ;
        RECT 1516.630 981.990 1517.810 983.170 ;
        RECT 1518.230 981.990 1519.410 983.170 ;
        RECT 1516.630 803.590 1517.810 804.770 ;
        RECT 1518.230 803.590 1519.410 804.770 ;
        RECT 1516.630 801.990 1517.810 803.170 ;
        RECT 1518.230 801.990 1519.410 803.170 ;
        RECT 1516.630 623.590 1517.810 624.770 ;
        RECT 1518.230 623.590 1519.410 624.770 ;
        RECT 1516.630 621.990 1517.810 623.170 ;
        RECT 1518.230 621.990 1519.410 623.170 ;
        RECT 1516.630 443.590 1517.810 444.770 ;
        RECT 1518.230 443.590 1519.410 444.770 ;
        RECT 1516.630 441.990 1517.810 443.170 ;
        RECT 1518.230 441.990 1519.410 443.170 ;
        RECT 1516.630 263.590 1517.810 264.770 ;
        RECT 1518.230 263.590 1519.410 264.770 ;
        RECT 1516.630 261.990 1517.810 263.170 ;
        RECT 1518.230 261.990 1519.410 263.170 ;
        RECT 1516.630 83.590 1517.810 84.770 ;
        RECT 1518.230 83.590 1519.410 84.770 ;
        RECT 1516.630 81.990 1517.810 83.170 ;
        RECT 1518.230 81.990 1519.410 83.170 ;
        RECT 1516.630 -17.310 1517.810 -16.130 ;
        RECT 1518.230 -17.310 1519.410 -16.130 ;
        RECT 1516.630 -18.910 1517.810 -17.730 ;
        RECT 1518.230 -18.910 1519.410 -17.730 ;
        RECT 1696.630 3537.410 1697.810 3538.590 ;
        RECT 1698.230 3537.410 1699.410 3538.590 ;
        RECT 1696.630 3535.810 1697.810 3536.990 ;
        RECT 1698.230 3535.810 1699.410 3536.990 ;
        RECT 1696.630 3503.590 1697.810 3504.770 ;
        RECT 1698.230 3503.590 1699.410 3504.770 ;
        RECT 1696.630 3501.990 1697.810 3503.170 ;
        RECT 1698.230 3501.990 1699.410 3503.170 ;
        RECT 1696.630 3323.590 1697.810 3324.770 ;
        RECT 1698.230 3323.590 1699.410 3324.770 ;
        RECT 1696.630 3321.990 1697.810 3323.170 ;
        RECT 1698.230 3321.990 1699.410 3323.170 ;
        RECT 1696.630 3143.590 1697.810 3144.770 ;
        RECT 1698.230 3143.590 1699.410 3144.770 ;
        RECT 1696.630 3141.990 1697.810 3143.170 ;
        RECT 1698.230 3141.990 1699.410 3143.170 ;
        RECT 1696.630 2963.590 1697.810 2964.770 ;
        RECT 1698.230 2963.590 1699.410 2964.770 ;
        RECT 1696.630 2961.990 1697.810 2963.170 ;
        RECT 1698.230 2961.990 1699.410 2963.170 ;
        RECT 1696.630 2783.590 1697.810 2784.770 ;
        RECT 1698.230 2783.590 1699.410 2784.770 ;
        RECT 1696.630 2781.990 1697.810 2783.170 ;
        RECT 1698.230 2781.990 1699.410 2783.170 ;
        RECT 1696.630 2603.590 1697.810 2604.770 ;
        RECT 1698.230 2603.590 1699.410 2604.770 ;
        RECT 1696.630 2601.990 1697.810 2603.170 ;
        RECT 1698.230 2601.990 1699.410 2603.170 ;
        RECT 1696.630 2423.590 1697.810 2424.770 ;
        RECT 1698.230 2423.590 1699.410 2424.770 ;
        RECT 1696.630 2421.990 1697.810 2423.170 ;
        RECT 1698.230 2421.990 1699.410 2423.170 ;
        RECT 1696.630 2243.590 1697.810 2244.770 ;
        RECT 1698.230 2243.590 1699.410 2244.770 ;
        RECT 1696.630 2241.990 1697.810 2243.170 ;
        RECT 1698.230 2241.990 1699.410 2243.170 ;
        RECT 1696.630 2063.590 1697.810 2064.770 ;
        RECT 1698.230 2063.590 1699.410 2064.770 ;
        RECT 1696.630 2061.990 1697.810 2063.170 ;
        RECT 1698.230 2061.990 1699.410 2063.170 ;
        RECT 1696.630 1883.590 1697.810 1884.770 ;
        RECT 1698.230 1883.590 1699.410 1884.770 ;
        RECT 1696.630 1881.990 1697.810 1883.170 ;
        RECT 1698.230 1881.990 1699.410 1883.170 ;
        RECT 1696.630 1703.590 1697.810 1704.770 ;
        RECT 1698.230 1703.590 1699.410 1704.770 ;
        RECT 1696.630 1701.990 1697.810 1703.170 ;
        RECT 1698.230 1701.990 1699.410 1703.170 ;
        RECT 1696.630 1523.590 1697.810 1524.770 ;
        RECT 1698.230 1523.590 1699.410 1524.770 ;
        RECT 1696.630 1521.990 1697.810 1523.170 ;
        RECT 1698.230 1521.990 1699.410 1523.170 ;
        RECT 1696.630 1343.590 1697.810 1344.770 ;
        RECT 1698.230 1343.590 1699.410 1344.770 ;
        RECT 1696.630 1341.990 1697.810 1343.170 ;
        RECT 1698.230 1341.990 1699.410 1343.170 ;
        RECT 1696.630 1163.590 1697.810 1164.770 ;
        RECT 1698.230 1163.590 1699.410 1164.770 ;
        RECT 1696.630 1161.990 1697.810 1163.170 ;
        RECT 1698.230 1161.990 1699.410 1163.170 ;
        RECT 1696.630 983.590 1697.810 984.770 ;
        RECT 1698.230 983.590 1699.410 984.770 ;
        RECT 1696.630 981.990 1697.810 983.170 ;
        RECT 1698.230 981.990 1699.410 983.170 ;
        RECT 1696.630 803.590 1697.810 804.770 ;
        RECT 1698.230 803.590 1699.410 804.770 ;
        RECT 1696.630 801.990 1697.810 803.170 ;
        RECT 1698.230 801.990 1699.410 803.170 ;
        RECT 1696.630 623.590 1697.810 624.770 ;
        RECT 1698.230 623.590 1699.410 624.770 ;
        RECT 1696.630 621.990 1697.810 623.170 ;
        RECT 1698.230 621.990 1699.410 623.170 ;
        RECT 1696.630 443.590 1697.810 444.770 ;
        RECT 1698.230 443.590 1699.410 444.770 ;
        RECT 1696.630 441.990 1697.810 443.170 ;
        RECT 1698.230 441.990 1699.410 443.170 ;
        RECT 1696.630 263.590 1697.810 264.770 ;
        RECT 1698.230 263.590 1699.410 264.770 ;
        RECT 1696.630 261.990 1697.810 263.170 ;
        RECT 1698.230 261.990 1699.410 263.170 ;
        RECT 1696.630 83.590 1697.810 84.770 ;
        RECT 1698.230 83.590 1699.410 84.770 ;
        RECT 1696.630 81.990 1697.810 83.170 ;
        RECT 1698.230 81.990 1699.410 83.170 ;
        RECT 1696.630 -17.310 1697.810 -16.130 ;
        RECT 1698.230 -17.310 1699.410 -16.130 ;
        RECT 1696.630 -18.910 1697.810 -17.730 ;
        RECT 1698.230 -18.910 1699.410 -17.730 ;
        RECT 1876.630 3537.410 1877.810 3538.590 ;
        RECT 1878.230 3537.410 1879.410 3538.590 ;
        RECT 1876.630 3535.810 1877.810 3536.990 ;
        RECT 1878.230 3535.810 1879.410 3536.990 ;
        RECT 1876.630 3503.590 1877.810 3504.770 ;
        RECT 1878.230 3503.590 1879.410 3504.770 ;
        RECT 1876.630 3501.990 1877.810 3503.170 ;
        RECT 1878.230 3501.990 1879.410 3503.170 ;
        RECT 1876.630 3323.590 1877.810 3324.770 ;
        RECT 1878.230 3323.590 1879.410 3324.770 ;
        RECT 1876.630 3321.990 1877.810 3323.170 ;
        RECT 1878.230 3321.990 1879.410 3323.170 ;
        RECT 1876.630 3143.590 1877.810 3144.770 ;
        RECT 1878.230 3143.590 1879.410 3144.770 ;
        RECT 1876.630 3141.990 1877.810 3143.170 ;
        RECT 1878.230 3141.990 1879.410 3143.170 ;
        RECT 1876.630 2963.590 1877.810 2964.770 ;
        RECT 1878.230 2963.590 1879.410 2964.770 ;
        RECT 1876.630 2961.990 1877.810 2963.170 ;
        RECT 1878.230 2961.990 1879.410 2963.170 ;
        RECT 1876.630 2783.590 1877.810 2784.770 ;
        RECT 1878.230 2783.590 1879.410 2784.770 ;
        RECT 1876.630 2781.990 1877.810 2783.170 ;
        RECT 1878.230 2781.990 1879.410 2783.170 ;
        RECT 1876.630 2603.590 1877.810 2604.770 ;
        RECT 1878.230 2603.590 1879.410 2604.770 ;
        RECT 1876.630 2601.990 1877.810 2603.170 ;
        RECT 1878.230 2601.990 1879.410 2603.170 ;
        RECT 1876.630 2423.590 1877.810 2424.770 ;
        RECT 1878.230 2423.590 1879.410 2424.770 ;
        RECT 1876.630 2421.990 1877.810 2423.170 ;
        RECT 1878.230 2421.990 1879.410 2423.170 ;
        RECT 1876.630 2243.590 1877.810 2244.770 ;
        RECT 1878.230 2243.590 1879.410 2244.770 ;
        RECT 1876.630 2241.990 1877.810 2243.170 ;
        RECT 1878.230 2241.990 1879.410 2243.170 ;
        RECT 1876.630 2063.590 1877.810 2064.770 ;
        RECT 1878.230 2063.590 1879.410 2064.770 ;
        RECT 1876.630 2061.990 1877.810 2063.170 ;
        RECT 1878.230 2061.990 1879.410 2063.170 ;
        RECT 1876.630 1883.590 1877.810 1884.770 ;
        RECT 1878.230 1883.590 1879.410 1884.770 ;
        RECT 1876.630 1881.990 1877.810 1883.170 ;
        RECT 1878.230 1881.990 1879.410 1883.170 ;
        RECT 1876.630 1703.590 1877.810 1704.770 ;
        RECT 1878.230 1703.590 1879.410 1704.770 ;
        RECT 1876.630 1701.990 1877.810 1703.170 ;
        RECT 1878.230 1701.990 1879.410 1703.170 ;
        RECT 1876.630 1523.590 1877.810 1524.770 ;
        RECT 1878.230 1523.590 1879.410 1524.770 ;
        RECT 1876.630 1521.990 1877.810 1523.170 ;
        RECT 1878.230 1521.990 1879.410 1523.170 ;
        RECT 1876.630 1343.590 1877.810 1344.770 ;
        RECT 1878.230 1343.590 1879.410 1344.770 ;
        RECT 1876.630 1341.990 1877.810 1343.170 ;
        RECT 1878.230 1341.990 1879.410 1343.170 ;
        RECT 1876.630 1163.590 1877.810 1164.770 ;
        RECT 1878.230 1163.590 1879.410 1164.770 ;
        RECT 1876.630 1161.990 1877.810 1163.170 ;
        RECT 1878.230 1161.990 1879.410 1163.170 ;
        RECT 1876.630 983.590 1877.810 984.770 ;
        RECT 1878.230 983.590 1879.410 984.770 ;
        RECT 1876.630 981.990 1877.810 983.170 ;
        RECT 1878.230 981.990 1879.410 983.170 ;
        RECT 1876.630 803.590 1877.810 804.770 ;
        RECT 1878.230 803.590 1879.410 804.770 ;
        RECT 1876.630 801.990 1877.810 803.170 ;
        RECT 1878.230 801.990 1879.410 803.170 ;
        RECT 1876.630 623.590 1877.810 624.770 ;
        RECT 1878.230 623.590 1879.410 624.770 ;
        RECT 1876.630 621.990 1877.810 623.170 ;
        RECT 1878.230 621.990 1879.410 623.170 ;
        RECT 1876.630 443.590 1877.810 444.770 ;
        RECT 1878.230 443.590 1879.410 444.770 ;
        RECT 1876.630 441.990 1877.810 443.170 ;
        RECT 1878.230 441.990 1879.410 443.170 ;
        RECT 1876.630 263.590 1877.810 264.770 ;
        RECT 1878.230 263.590 1879.410 264.770 ;
        RECT 1876.630 261.990 1877.810 263.170 ;
        RECT 1878.230 261.990 1879.410 263.170 ;
        RECT 1876.630 83.590 1877.810 84.770 ;
        RECT 1878.230 83.590 1879.410 84.770 ;
        RECT 1876.630 81.990 1877.810 83.170 ;
        RECT 1878.230 81.990 1879.410 83.170 ;
        RECT 1876.630 -17.310 1877.810 -16.130 ;
        RECT 1878.230 -17.310 1879.410 -16.130 ;
        RECT 1876.630 -18.910 1877.810 -17.730 ;
        RECT 1878.230 -18.910 1879.410 -17.730 ;
        RECT 2056.630 3537.410 2057.810 3538.590 ;
        RECT 2058.230 3537.410 2059.410 3538.590 ;
        RECT 2056.630 3535.810 2057.810 3536.990 ;
        RECT 2058.230 3535.810 2059.410 3536.990 ;
        RECT 2056.630 3503.590 2057.810 3504.770 ;
        RECT 2058.230 3503.590 2059.410 3504.770 ;
        RECT 2056.630 3501.990 2057.810 3503.170 ;
        RECT 2058.230 3501.990 2059.410 3503.170 ;
        RECT 2056.630 3323.590 2057.810 3324.770 ;
        RECT 2058.230 3323.590 2059.410 3324.770 ;
        RECT 2056.630 3321.990 2057.810 3323.170 ;
        RECT 2058.230 3321.990 2059.410 3323.170 ;
        RECT 2056.630 3143.590 2057.810 3144.770 ;
        RECT 2058.230 3143.590 2059.410 3144.770 ;
        RECT 2056.630 3141.990 2057.810 3143.170 ;
        RECT 2058.230 3141.990 2059.410 3143.170 ;
        RECT 2056.630 2963.590 2057.810 2964.770 ;
        RECT 2058.230 2963.590 2059.410 2964.770 ;
        RECT 2056.630 2961.990 2057.810 2963.170 ;
        RECT 2058.230 2961.990 2059.410 2963.170 ;
        RECT 2056.630 2783.590 2057.810 2784.770 ;
        RECT 2058.230 2783.590 2059.410 2784.770 ;
        RECT 2056.630 2781.990 2057.810 2783.170 ;
        RECT 2058.230 2781.990 2059.410 2783.170 ;
        RECT 2056.630 2603.590 2057.810 2604.770 ;
        RECT 2058.230 2603.590 2059.410 2604.770 ;
        RECT 2056.630 2601.990 2057.810 2603.170 ;
        RECT 2058.230 2601.990 2059.410 2603.170 ;
        RECT 2056.630 2423.590 2057.810 2424.770 ;
        RECT 2058.230 2423.590 2059.410 2424.770 ;
        RECT 2056.630 2421.990 2057.810 2423.170 ;
        RECT 2058.230 2421.990 2059.410 2423.170 ;
        RECT 2056.630 2243.590 2057.810 2244.770 ;
        RECT 2058.230 2243.590 2059.410 2244.770 ;
        RECT 2056.630 2241.990 2057.810 2243.170 ;
        RECT 2058.230 2241.990 2059.410 2243.170 ;
        RECT 2056.630 2063.590 2057.810 2064.770 ;
        RECT 2058.230 2063.590 2059.410 2064.770 ;
        RECT 2056.630 2061.990 2057.810 2063.170 ;
        RECT 2058.230 2061.990 2059.410 2063.170 ;
        RECT 2056.630 1883.590 2057.810 1884.770 ;
        RECT 2058.230 1883.590 2059.410 1884.770 ;
        RECT 2056.630 1881.990 2057.810 1883.170 ;
        RECT 2058.230 1881.990 2059.410 1883.170 ;
        RECT 2056.630 1703.590 2057.810 1704.770 ;
        RECT 2058.230 1703.590 2059.410 1704.770 ;
        RECT 2056.630 1701.990 2057.810 1703.170 ;
        RECT 2058.230 1701.990 2059.410 1703.170 ;
        RECT 2056.630 1523.590 2057.810 1524.770 ;
        RECT 2058.230 1523.590 2059.410 1524.770 ;
        RECT 2056.630 1521.990 2057.810 1523.170 ;
        RECT 2058.230 1521.990 2059.410 1523.170 ;
        RECT 2056.630 1343.590 2057.810 1344.770 ;
        RECT 2058.230 1343.590 2059.410 1344.770 ;
        RECT 2056.630 1341.990 2057.810 1343.170 ;
        RECT 2058.230 1341.990 2059.410 1343.170 ;
        RECT 2056.630 1163.590 2057.810 1164.770 ;
        RECT 2058.230 1163.590 2059.410 1164.770 ;
        RECT 2056.630 1161.990 2057.810 1163.170 ;
        RECT 2058.230 1161.990 2059.410 1163.170 ;
        RECT 2056.630 983.590 2057.810 984.770 ;
        RECT 2058.230 983.590 2059.410 984.770 ;
        RECT 2056.630 981.990 2057.810 983.170 ;
        RECT 2058.230 981.990 2059.410 983.170 ;
        RECT 2056.630 803.590 2057.810 804.770 ;
        RECT 2058.230 803.590 2059.410 804.770 ;
        RECT 2056.630 801.990 2057.810 803.170 ;
        RECT 2058.230 801.990 2059.410 803.170 ;
        RECT 2056.630 623.590 2057.810 624.770 ;
        RECT 2058.230 623.590 2059.410 624.770 ;
        RECT 2056.630 621.990 2057.810 623.170 ;
        RECT 2058.230 621.990 2059.410 623.170 ;
        RECT 2056.630 443.590 2057.810 444.770 ;
        RECT 2058.230 443.590 2059.410 444.770 ;
        RECT 2056.630 441.990 2057.810 443.170 ;
        RECT 2058.230 441.990 2059.410 443.170 ;
        RECT 2056.630 263.590 2057.810 264.770 ;
        RECT 2058.230 263.590 2059.410 264.770 ;
        RECT 2056.630 261.990 2057.810 263.170 ;
        RECT 2058.230 261.990 2059.410 263.170 ;
        RECT 2056.630 83.590 2057.810 84.770 ;
        RECT 2058.230 83.590 2059.410 84.770 ;
        RECT 2056.630 81.990 2057.810 83.170 ;
        RECT 2058.230 81.990 2059.410 83.170 ;
        RECT 2056.630 -17.310 2057.810 -16.130 ;
        RECT 2058.230 -17.310 2059.410 -16.130 ;
        RECT 2056.630 -18.910 2057.810 -17.730 ;
        RECT 2058.230 -18.910 2059.410 -17.730 ;
        RECT 2236.630 3537.410 2237.810 3538.590 ;
        RECT 2238.230 3537.410 2239.410 3538.590 ;
        RECT 2236.630 3535.810 2237.810 3536.990 ;
        RECT 2238.230 3535.810 2239.410 3536.990 ;
        RECT 2236.630 3503.590 2237.810 3504.770 ;
        RECT 2238.230 3503.590 2239.410 3504.770 ;
        RECT 2236.630 3501.990 2237.810 3503.170 ;
        RECT 2238.230 3501.990 2239.410 3503.170 ;
        RECT 2236.630 3323.590 2237.810 3324.770 ;
        RECT 2238.230 3323.590 2239.410 3324.770 ;
        RECT 2236.630 3321.990 2237.810 3323.170 ;
        RECT 2238.230 3321.990 2239.410 3323.170 ;
        RECT 2236.630 3143.590 2237.810 3144.770 ;
        RECT 2238.230 3143.590 2239.410 3144.770 ;
        RECT 2236.630 3141.990 2237.810 3143.170 ;
        RECT 2238.230 3141.990 2239.410 3143.170 ;
        RECT 2236.630 2963.590 2237.810 2964.770 ;
        RECT 2238.230 2963.590 2239.410 2964.770 ;
        RECT 2236.630 2961.990 2237.810 2963.170 ;
        RECT 2238.230 2961.990 2239.410 2963.170 ;
        RECT 2236.630 2783.590 2237.810 2784.770 ;
        RECT 2238.230 2783.590 2239.410 2784.770 ;
        RECT 2236.630 2781.990 2237.810 2783.170 ;
        RECT 2238.230 2781.990 2239.410 2783.170 ;
        RECT 2236.630 2603.590 2237.810 2604.770 ;
        RECT 2238.230 2603.590 2239.410 2604.770 ;
        RECT 2236.630 2601.990 2237.810 2603.170 ;
        RECT 2238.230 2601.990 2239.410 2603.170 ;
        RECT 2236.630 2423.590 2237.810 2424.770 ;
        RECT 2238.230 2423.590 2239.410 2424.770 ;
        RECT 2236.630 2421.990 2237.810 2423.170 ;
        RECT 2238.230 2421.990 2239.410 2423.170 ;
        RECT 2236.630 2243.590 2237.810 2244.770 ;
        RECT 2238.230 2243.590 2239.410 2244.770 ;
        RECT 2236.630 2241.990 2237.810 2243.170 ;
        RECT 2238.230 2241.990 2239.410 2243.170 ;
        RECT 2236.630 2063.590 2237.810 2064.770 ;
        RECT 2238.230 2063.590 2239.410 2064.770 ;
        RECT 2236.630 2061.990 2237.810 2063.170 ;
        RECT 2238.230 2061.990 2239.410 2063.170 ;
        RECT 2236.630 1883.590 2237.810 1884.770 ;
        RECT 2238.230 1883.590 2239.410 1884.770 ;
        RECT 2236.630 1881.990 2237.810 1883.170 ;
        RECT 2238.230 1881.990 2239.410 1883.170 ;
        RECT 2236.630 1703.590 2237.810 1704.770 ;
        RECT 2238.230 1703.590 2239.410 1704.770 ;
        RECT 2236.630 1701.990 2237.810 1703.170 ;
        RECT 2238.230 1701.990 2239.410 1703.170 ;
        RECT 2236.630 1523.590 2237.810 1524.770 ;
        RECT 2238.230 1523.590 2239.410 1524.770 ;
        RECT 2236.630 1521.990 2237.810 1523.170 ;
        RECT 2238.230 1521.990 2239.410 1523.170 ;
        RECT 2236.630 1343.590 2237.810 1344.770 ;
        RECT 2238.230 1343.590 2239.410 1344.770 ;
        RECT 2236.630 1341.990 2237.810 1343.170 ;
        RECT 2238.230 1341.990 2239.410 1343.170 ;
        RECT 2236.630 1163.590 2237.810 1164.770 ;
        RECT 2238.230 1163.590 2239.410 1164.770 ;
        RECT 2236.630 1161.990 2237.810 1163.170 ;
        RECT 2238.230 1161.990 2239.410 1163.170 ;
        RECT 2236.630 983.590 2237.810 984.770 ;
        RECT 2238.230 983.590 2239.410 984.770 ;
        RECT 2236.630 981.990 2237.810 983.170 ;
        RECT 2238.230 981.990 2239.410 983.170 ;
        RECT 2236.630 803.590 2237.810 804.770 ;
        RECT 2238.230 803.590 2239.410 804.770 ;
        RECT 2236.630 801.990 2237.810 803.170 ;
        RECT 2238.230 801.990 2239.410 803.170 ;
        RECT 2236.630 623.590 2237.810 624.770 ;
        RECT 2238.230 623.590 2239.410 624.770 ;
        RECT 2236.630 621.990 2237.810 623.170 ;
        RECT 2238.230 621.990 2239.410 623.170 ;
        RECT 2236.630 443.590 2237.810 444.770 ;
        RECT 2238.230 443.590 2239.410 444.770 ;
        RECT 2236.630 441.990 2237.810 443.170 ;
        RECT 2238.230 441.990 2239.410 443.170 ;
        RECT 2236.630 263.590 2237.810 264.770 ;
        RECT 2238.230 263.590 2239.410 264.770 ;
        RECT 2236.630 261.990 2237.810 263.170 ;
        RECT 2238.230 261.990 2239.410 263.170 ;
        RECT 2236.630 83.590 2237.810 84.770 ;
        RECT 2238.230 83.590 2239.410 84.770 ;
        RECT 2236.630 81.990 2237.810 83.170 ;
        RECT 2238.230 81.990 2239.410 83.170 ;
        RECT 2236.630 -17.310 2237.810 -16.130 ;
        RECT 2238.230 -17.310 2239.410 -16.130 ;
        RECT 2236.630 -18.910 2237.810 -17.730 ;
        RECT 2238.230 -18.910 2239.410 -17.730 ;
        RECT 2416.630 3537.410 2417.810 3538.590 ;
        RECT 2418.230 3537.410 2419.410 3538.590 ;
        RECT 2416.630 3535.810 2417.810 3536.990 ;
        RECT 2418.230 3535.810 2419.410 3536.990 ;
        RECT 2416.630 3503.590 2417.810 3504.770 ;
        RECT 2418.230 3503.590 2419.410 3504.770 ;
        RECT 2416.630 3501.990 2417.810 3503.170 ;
        RECT 2418.230 3501.990 2419.410 3503.170 ;
        RECT 2416.630 3323.590 2417.810 3324.770 ;
        RECT 2418.230 3323.590 2419.410 3324.770 ;
        RECT 2416.630 3321.990 2417.810 3323.170 ;
        RECT 2418.230 3321.990 2419.410 3323.170 ;
        RECT 2416.630 3143.590 2417.810 3144.770 ;
        RECT 2418.230 3143.590 2419.410 3144.770 ;
        RECT 2416.630 3141.990 2417.810 3143.170 ;
        RECT 2418.230 3141.990 2419.410 3143.170 ;
        RECT 2416.630 2963.590 2417.810 2964.770 ;
        RECT 2418.230 2963.590 2419.410 2964.770 ;
        RECT 2416.630 2961.990 2417.810 2963.170 ;
        RECT 2418.230 2961.990 2419.410 2963.170 ;
        RECT 2416.630 2783.590 2417.810 2784.770 ;
        RECT 2418.230 2783.590 2419.410 2784.770 ;
        RECT 2416.630 2781.990 2417.810 2783.170 ;
        RECT 2418.230 2781.990 2419.410 2783.170 ;
        RECT 2416.630 2603.590 2417.810 2604.770 ;
        RECT 2418.230 2603.590 2419.410 2604.770 ;
        RECT 2416.630 2601.990 2417.810 2603.170 ;
        RECT 2418.230 2601.990 2419.410 2603.170 ;
        RECT 2416.630 2423.590 2417.810 2424.770 ;
        RECT 2418.230 2423.590 2419.410 2424.770 ;
        RECT 2416.630 2421.990 2417.810 2423.170 ;
        RECT 2418.230 2421.990 2419.410 2423.170 ;
        RECT 2416.630 2243.590 2417.810 2244.770 ;
        RECT 2418.230 2243.590 2419.410 2244.770 ;
        RECT 2416.630 2241.990 2417.810 2243.170 ;
        RECT 2418.230 2241.990 2419.410 2243.170 ;
        RECT 2416.630 2063.590 2417.810 2064.770 ;
        RECT 2418.230 2063.590 2419.410 2064.770 ;
        RECT 2416.630 2061.990 2417.810 2063.170 ;
        RECT 2418.230 2061.990 2419.410 2063.170 ;
        RECT 2416.630 1883.590 2417.810 1884.770 ;
        RECT 2418.230 1883.590 2419.410 1884.770 ;
        RECT 2416.630 1881.990 2417.810 1883.170 ;
        RECT 2418.230 1881.990 2419.410 1883.170 ;
        RECT 2416.630 1703.590 2417.810 1704.770 ;
        RECT 2418.230 1703.590 2419.410 1704.770 ;
        RECT 2416.630 1701.990 2417.810 1703.170 ;
        RECT 2418.230 1701.990 2419.410 1703.170 ;
        RECT 2416.630 1523.590 2417.810 1524.770 ;
        RECT 2418.230 1523.590 2419.410 1524.770 ;
        RECT 2416.630 1521.990 2417.810 1523.170 ;
        RECT 2418.230 1521.990 2419.410 1523.170 ;
        RECT 2416.630 1343.590 2417.810 1344.770 ;
        RECT 2418.230 1343.590 2419.410 1344.770 ;
        RECT 2416.630 1341.990 2417.810 1343.170 ;
        RECT 2418.230 1341.990 2419.410 1343.170 ;
        RECT 2416.630 1163.590 2417.810 1164.770 ;
        RECT 2418.230 1163.590 2419.410 1164.770 ;
        RECT 2416.630 1161.990 2417.810 1163.170 ;
        RECT 2418.230 1161.990 2419.410 1163.170 ;
        RECT 2416.630 983.590 2417.810 984.770 ;
        RECT 2418.230 983.590 2419.410 984.770 ;
        RECT 2416.630 981.990 2417.810 983.170 ;
        RECT 2418.230 981.990 2419.410 983.170 ;
        RECT 2416.630 803.590 2417.810 804.770 ;
        RECT 2418.230 803.590 2419.410 804.770 ;
        RECT 2416.630 801.990 2417.810 803.170 ;
        RECT 2418.230 801.990 2419.410 803.170 ;
        RECT 2416.630 623.590 2417.810 624.770 ;
        RECT 2418.230 623.590 2419.410 624.770 ;
        RECT 2416.630 621.990 2417.810 623.170 ;
        RECT 2418.230 621.990 2419.410 623.170 ;
        RECT 2416.630 443.590 2417.810 444.770 ;
        RECT 2418.230 443.590 2419.410 444.770 ;
        RECT 2416.630 441.990 2417.810 443.170 ;
        RECT 2418.230 441.990 2419.410 443.170 ;
        RECT 2416.630 263.590 2417.810 264.770 ;
        RECT 2418.230 263.590 2419.410 264.770 ;
        RECT 2416.630 261.990 2417.810 263.170 ;
        RECT 2418.230 261.990 2419.410 263.170 ;
        RECT 2416.630 83.590 2417.810 84.770 ;
        RECT 2418.230 83.590 2419.410 84.770 ;
        RECT 2416.630 81.990 2417.810 83.170 ;
        RECT 2418.230 81.990 2419.410 83.170 ;
        RECT 2416.630 -17.310 2417.810 -16.130 ;
        RECT 2418.230 -17.310 2419.410 -16.130 ;
        RECT 2416.630 -18.910 2417.810 -17.730 ;
        RECT 2418.230 -18.910 2419.410 -17.730 ;
        RECT 2596.630 3537.410 2597.810 3538.590 ;
        RECT 2598.230 3537.410 2599.410 3538.590 ;
        RECT 2596.630 3535.810 2597.810 3536.990 ;
        RECT 2598.230 3535.810 2599.410 3536.990 ;
        RECT 2596.630 3503.590 2597.810 3504.770 ;
        RECT 2598.230 3503.590 2599.410 3504.770 ;
        RECT 2596.630 3501.990 2597.810 3503.170 ;
        RECT 2598.230 3501.990 2599.410 3503.170 ;
        RECT 2596.630 3323.590 2597.810 3324.770 ;
        RECT 2598.230 3323.590 2599.410 3324.770 ;
        RECT 2596.630 3321.990 2597.810 3323.170 ;
        RECT 2598.230 3321.990 2599.410 3323.170 ;
        RECT 2596.630 3143.590 2597.810 3144.770 ;
        RECT 2598.230 3143.590 2599.410 3144.770 ;
        RECT 2596.630 3141.990 2597.810 3143.170 ;
        RECT 2598.230 3141.990 2599.410 3143.170 ;
        RECT 2596.630 2963.590 2597.810 2964.770 ;
        RECT 2598.230 2963.590 2599.410 2964.770 ;
        RECT 2596.630 2961.990 2597.810 2963.170 ;
        RECT 2598.230 2961.990 2599.410 2963.170 ;
        RECT 2596.630 2783.590 2597.810 2784.770 ;
        RECT 2598.230 2783.590 2599.410 2784.770 ;
        RECT 2596.630 2781.990 2597.810 2783.170 ;
        RECT 2598.230 2781.990 2599.410 2783.170 ;
        RECT 2596.630 2603.590 2597.810 2604.770 ;
        RECT 2598.230 2603.590 2599.410 2604.770 ;
        RECT 2596.630 2601.990 2597.810 2603.170 ;
        RECT 2598.230 2601.990 2599.410 2603.170 ;
        RECT 2596.630 2423.590 2597.810 2424.770 ;
        RECT 2598.230 2423.590 2599.410 2424.770 ;
        RECT 2596.630 2421.990 2597.810 2423.170 ;
        RECT 2598.230 2421.990 2599.410 2423.170 ;
        RECT 2596.630 2243.590 2597.810 2244.770 ;
        RECT 2598.230 2243.590 2599.410 2244.770 ;
        RECT 2596.630 2241.990 2597.810 2243.170 ;
        RECT 2598.230 2241.990 2599.410 2243.170 ;
        RECT 2596.630 2063.590 2597.810 2064.770 ;
        RECT 2598.230 2063.590 2599.410 2064.770 ;
        RECT 2596.630 2061.990 2597.810 2063.170 ;
        RECT 2598.230 2061.990 2599.410 2063.170 ;
        RECT 2596.630 1883.590 2597.810 1884.770 ;
        RECT 2598.230 1883.590 2599.410 1884.770 ;
        RECT 2596.630 1881.990 2597.810 1883.170 ;
        RECT 2598.230 1881.990 2599.410 1883.170 ;
        RECT 2596.630 1703.590 2597.810 1704.770 ;
        RECT 2598.230 1703.590 2599.410 1704.770 ;
        RECT 2596.630 1701.990 2597.810 1703.170 ;
        RECT 2598.230 1701.990 2599.410 1703.170 ;
        RECT 2596.630 1523.590 2597.810 1524.770 ;
        RECT 2598.230 1523.590 2599.410 1524.770 ;
        RECT 2596.630 1521.990 2597.810 1523.170 ;
        RECT 2598.230 1521.990 2599.410 1523.170 ;
        RECT 2596.630 1343.590 2597.810 1344.770 ;
        RECT 2598.230 1343.590 2599.410 1344.770 ;
        RECT 2596.630 1341.990 2597.810 1343.170 ;
        RECT 2598.230 1341.990 2599.410 1343.170 ;
        RECT 2596.630 1163.590 2597.810 1164.770 ;
        RECT 2598.230 1163.590 2599.410 1164.770 ;
        RECT 2596.630 1161.990 2597.810 1163.170 ;
        RECT 2598.230 1161.990 2599.410 1163.170 ;
        RECT 2596.630 983.590 2597.810 984.770 ;
        RECT 2598.230 983.590 2599.410 984.770 ;
        RECT 2596.630 981.990 2597.810 983.170 ;
        RECT 2598.230 981.990 2599.410 983.170 ;
        RECT 2596.630 803.590 2597.810 804.770 ;
        RECT 2598.230 803.590 2599.410 804.770 ;
        RECT 2596.630 801.990 2597.810 803.170 ;
        RECT 2598.230 801.990 2599.410 803.170 ;
        RECT 2596.630 623.590 2597.810 624.770 ;
        RECT 2598.230 623.590 2599.410 624.770 ;
        RECT 2596.630 621.990 2597.810 623.170 ;
        RECT 2598.230 621.990 2599.410 623.170 ;
        RECT 2596.630 443.590 2597.810 444.770 ;
        RECT 2598.230 443.590 2599.410 444.770 ;
        RECT 2596.630 441.990 2597.810 443.170 ;
        RECT 2598.230 441.990 2599.410 443.170 ;
        RECT 2596.630 263.590 2597.810 264.770 ;
        RECT 2598.230 263.590 2599.410 264.770 ;
        RECT 2596.630 261.990 2597.810 263.170 ;
        RECT 2598.230 261.990 2599.410 263.170 ;
        RECT 2596.630 83.590 2597.810 84.770 ;
        RECT 2598.230 83.590 2599.410 84.770 ;
        RECT 2596.630 81.990 2597.810 83.170 ;
        RECT 2598.230 81.990 2599.410 83.170 ;
        RECT 2596.630 -17.310 2597.810 -16.130 ;
        RECT 2598.230 -17.310 2599.410 -16.130 ;
        RECT 2596.630 -18.910 2597.810 -17.730 ;
        RECT 2598.230 -18.910 2599.410 -17.730 ;
        RECT 2776.630 3537.410 2777.810 3538.590 ;
        RECT 2778.230 3537.410 2779.410 3538.590 ;
        RECT 2776.630 3535.810 2777.810 3536.990 ;
        RECT 2778.230 3535.810 2779.410 3536.990 ;
        RECT 2776.630 3503.590 2777.810 3504.770 ;
        RECT 2778.230 3503.590 2779.410 3504.770 ;
        RECT 2776.630 3501.990 2777.810 3503.170 ;
        RECT 2778.230 3501.990 2779.410 3503.170 ;
        RECT 2776.630 3323.590 2777.810 3324.770 ;
        RECT 2778.230 3323.590 2779.410 3324.770 ;
        RECT 2776.630 3321.990 2777.810 3323.170 ;
        RECT 2778.230 3321.990 2779.410 3323.170 ;
        RECT 2776.630 3143.590 2777.810 3144.770 ;
        RECT 2778.230 3143.590 2779.410 3144.770 ;
        RECT 2776.630 3141.990 2777.810 3143.170 ;
        RECT 2778.230 3141.990 2779.410 3143.170 ;
        RECT 2776.630 2963.590 2777.810 2964.770 ;
        RECT 2778.230 2963.590 2779.410 2964.770 ;
        RECT 2776.630 2961.990 2777.810 2963.170 ;
        RECT 2778.230 2961.990 2779.410 2963.170 ;
        RECT 2776.630 2783.590 2777.810 2784.770 ;
        RECT 2778.230 2783.590 2779.410 2784.770 ;
        RECT 2776.630 2781.990 2777.810 2783.170 ;
        RECT 2778.230 2781.990 2779.410 2783.170 ;
        RECT 2776.630 2603.590 2777.810 2604.770 ;
        RECT 2778.230 2603.590 2779.410 2604.770 ;
        RECT 2776.630 2601.990 2777.810 2603.170 ;
        RECT 2778.230 2601.990 2779.410 2603.170 ;
        RECT 2776.630 2423.590 2777.810 2424.770 ;
        RECT 2778.230 2423.590 2779.410 2424.770 ;
        RECT 2776.630 2421.990 2777.810 2423.170 ;
        RECT 2778.230 2421.990 2779.410 2423.170 ;
        RECT 2776.630 2243.590 2777.810 2244.770 ;
        RECT 2778.230 2243.590 2779.410 2244.770 ;
        RECT 2776.630 2241.990 2777.810 2243.170 ;
        RECT 2778.230 2241.990 2779.410 2243.170 ;
        RECT 2776.630 2063.590 2777.810 2064.770 ;
        RECT 2778.230 2063.590 2779.410 2064.770 ;
        RECT 2776.630 2061.990 2777.810 2063.170 ;
        RECT 2778.230 2061.990 2779.410 2063.170 ;
        RECT 2776.630 1883.590 2777.810 1884.770 ;
        RECT 2778.230 1883.590 2779.410 1884.770 ;
        RECT 2776.630 1881.990 2777.810 1883.170 ;
        RECT 2778.230 1881.990 2779.410 1883.170 ;
        RECT 2776.630 1703.590 2777.810 1704.770 ;
        RECT 2778.230 1703.590 2779.410 1704.770 ;
        RECT 2776.630 1701.990 2777.810 1703.170 ;
        RECT 2778.230 1701.990 2779.410 1703.170 ;
        RECT 2776.630 1523.590 2777.810 1524.770 ;
        RECT 2778.230 1523.590 2779.410 1524.770 ;
        RECT 2776.630 1521.990 2777.810 1523.170 ;
        RECT 2778.230 1521.990 2779.410 1523.170 ;
        RECT 2776.630 1343.590 2777.810 1344.770 ;
        RECT 2778.230 1343.590 2779.410 1344.770 ;
        RECT 2776.630 1341.990 2777.810 1343.170 ;
        RECT 2778.230 1341.990 2779.410 1343.170 ;
        RECT 2776.630 1163.590 2777.810 1164.770 ;
        RECT 2778.230 1163.590 2779.410 1164.770 ;
        RECT 2776.630 1161.990 2777.810 1163.170 ;
        RECT 2778.230 1161.990 2779.410 1163.170 ;
        RECT 2776.630 983.590 2777.810 984.770 ;
        RECT 2778.230 983.590 2779.410 984.770 ;
        RECT 2776.630 981.990 2777.810 983.170 ;
        RECT 2778.230 981.990 2779.410 983.170 ;
        RECT 2776.630 803.590 2777.810 804.770 ;
        RECT 2778.230 803.590 2779.410 804.770 ;
        RECT 2776.630 801.990 2777.810 803.170 ;
        RECT 2778.230 801.990 2779.410 803.170 ;
        RECT 2776.630 623.590 2777.810 624.770 ;
        RECT 2778.230 623.590 2779.410 624.770 ;
        RECT 2776.630 621.990 2777.810 623.170 ;
        RECT 2778.230 621.990 2779.410 623.170 ;
        RECT 2776.630 443.590 2777.810 444.770 ;
        RECT 2778.230 443.590 2779.410 444.770 ;
        RECT 2776.630 441.990 2777.810 443.170 ;
        RECT 2778.230 441.990 2779.410 443.170 ;
        RECT 2776.630 263.590 2777.810 264.770 ;
        RECT 2778.230 263.590 2779.410 264.770 ;
        RECT 2776.630 261.990 2777.810 263.170 ;
        RECT 2778.230 261.990 2779.410 263.170 ;
        RECT 2776.630 83.590 2777.810 84.770 ;
        RECT 2778.230 83.590 2779.410 84.770 ;
        RECT 2776.630 81.990 2777.810 83.170 ;
        RECT 2778.230 81.990 2779.410 83.170 ;
        RECT 2776.630 -17.310 2777.810 -16.130 ;
        RECT 2778.230 -17.310 2779.410 -16.130 ;
        RECT 2776.630 -18.910 2777.810 -17.730 ;
        RECT 2778.230 -18.910 2779.410 -17.730 ;
        RECT 2941.110 3537.410 2942.290 3538.590 ;
        RECT 2942.710 3537.410 2943.890 3538.590 ;
        RECT 2941.110 3535.810 2942.290 3536.990 ;
        RECT 2942.710 3535.810 2943.890 3536.990 ;
        RECT 2941.110 3503.590 2942.290 3504.770 ;
        RECT 2942.710 3503.590 2943.890 3504.770 ;
        RECT 2941.110 3501.990 2942.290 3503.170 ;
        RECT 2942.710 3501.990 2943.890 3503.170 ;
        RECT 2941.110 3323.590 2942.290 3324.770 ;
        RECT 2942.710 3323.590 2943.890 3324.770 ;
        RECT 2941.110 3321.990 2942.290 3323.170 ;
        RECT 2942.710 3321.990 2943.890 3323.170 ;
        RECT 2941.110 3143.590 2942.290 3144.770 ;
        RECT 2942.710 3143.590 2943.890 3144.770 ;
        RECT 2941.110 3141.990 2942.290 3143.170 ;
        RECT 2942.710 3141.990 2943.890 3143.170 ;
        RECT 2941.110 2963.590 2942.290 2964.770 ;
        RECT 2942.710 2963.590 2943.890 2964.770 ;
        RECT 2941.110 2961.990 2942.290 2963.170 ;
        RECT 2942.710 2961.990 2943.890 2963.170 ;
        RECT 2941.110 2783.590 2942.290 2784.770 ;
        RECT 2942.710 2783.590 2943.890 2784.770 ;
        RECT 2941.110 2781.990 2942.290 2783.170 ;
        RECT 2942.710 2781.990 2943.890 2783.170 ;
        RECT 2941.110 2603.590 2942.290 2604.770 ;
        RECT 2942.710 2603.590 2943.890 2604.770 ;
        RECT 2941.110 2601.990 2942.290 2603.170 ;
        RECT 2942.710 2601.990 2943.890 2603.170 ;
        RECT 2941.110 2423.590 2942.290 2424.770 ;
        RECT 2942.710 2423.590 2943.890 2424.770 ;
        RECT 2941.110 2421.990 2942.290 2423.170 ;
        RECT 2942.710 2421.990 2943.890 2423.170 ;
        RECT 2941.110 2243.590 2942.290 2244.770 ;
        RECT 2942.710 2243.590 2943.890 2244.770 ;
        RECT 2941.110 2241.990 2942.290 2243.170 ;
        RECT 2942.710 2241.990 2943.890 2243.170 ;
        RECT 2941.110 2063.590 2942.290 2064.770 ;
        RECT 2942.710 2063.590 2943.890 2064.770 ;
        RECT 2941.110 2061.990 2942.290 2063.170 ;
        RECT 2942.710 2061.990 2943.890 2063.170 ;
        RECT 2941.110 1883.590 2942.290 1884.770 ;
        RECT 2942.710 1883.590 2943.890 1884.770 ;
        RECT 2941.110 1881.990 2942.290 1883.170 ;
        RECT 2942.710 1881.990 2943.890 1883.170 ;
        RECT 2941.110 1703.590 2942.290 1704.770 ;
        RECT 2942.710 1703.590 2943.890 1704.770 ;
        RECT 2941.110 1701.990 2942.290 1703.170 ;
        RECT 2942.710 1701.990 2943.890 1703.170 ;
        RECT 2941.110 1523.590 2942.290 1524.770 ;
        RECT 2942.710 1523.590 2943.890 1524.770 ;
        RECT 2941.110 1521.990 2942.290 1523.170 ;
        RECT 2942.710 1521.990 2943.890 1523.170 ;
        RECT 2941.110 1343.590 2942.290 1344.770 ;
        RECT 2942.710 1343.590 2943.890 1344.770 ;
        RECT 2941.110 1341.990 2942.290 1343.170 ;
        RECT 2942.710 1341.990 2943.890 1343.170 ;
        RECT 2941.110 1163.590 2942.290 1164.770 ;
        RECT 2942.710 1163.590 2943.890 1164.770 ;
        RECT 2941.110 1161.990 2942.290 1163.170 ;
        RECT 2942.710 1161.990 2943.890 1163.170 ;
        RECT 2941.110 983.590 2942.290 984.770 ;
        RECT 2942.710 983.590 2943.890 984.770 ;
        RECT 2941.110 981.990 2942.290 983.170 ;
        RECT 2942.710 981.990 2943.890 983.170 ;
        RECT 2941.110 803.590 2942.290 804.770 ;
        RECT 2942.710 803.590 2943.890 804.770 ;
        RECT 2941.110 801.990 2942.290 803.170 ;
        RECT 2942.710 801.990 2943.890 803.170 ;
        RECT 2941.110 623.590 2942.290 624.770 ;
        RECT 2942.710 623.590 2943.890 624.770 ;
        RECT 2941.110 621.990 2942.290 623.170 ;
        RECT 2942.710 621.990 2943.890 623.170 ;
        RECT 2941.110 443.590 2942.290 444.770 ;
        RECT 2942.710 443.590 2943.890 444.770 ;
        RECT 2941.110 441.990 2942.290 443.170 ;
        RECT 2942.710 441.990 2943.890 443.170 ;
        RECT 2941.110 263.590 2942.290 264.770 ;
        RECT 2942.710 263.590 2943.890 264.770 ;
        RECT 2941.110 261.990 2942.290 263.170 ;
        RECT 2942.710 261.990 2943.890 263.170 ;
        RECT 2941.110 83.590 2942.290 84.770 ;
        RECT 2942.710 83.590 2943.890 84.770 ;
        RECT 2941.110 81.990 2942.290 83.170 ;
        RECT 2942.710 81.990 2943.890 83.170 ;
        RECT 2941.110 -17.310 2942.290 -16.130 ;
        RECT 2942.710 -17.310 2943.890 -16.130 ;
        RECT 2941.110 -18.910 2942.290 -17.730 ;
        RECT 2942.710 -18.910 2943.890 -17.730 ;
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
        RECT -43.630 3501.830 2963.250 3504.930 ;
        RECT -43.630 3321.830 2963.250 3324.930 ;
        RECT -43.630 3141.830 2963.250 3144.930 ;
        RECT -43.630 2961.830 2963.250 2964.930 ;
        RECT -43.630 2781.830 2963.250 2784.930 ;
        RECT -43.630 2601.830 2963.250 2604.930 ;
        RECT -43.630 2421.830 2963.250 2424.930 ;
        RECT -43.630 2241.830 2963.250 2244.930 ;
        RECT -43.630 2061.830 2963.250 2064.930 ;
        RECT -43.630 1881.830 2963.250 1884.930 ;
        RECT -43.630 1701.830 2963.250 1704.930 ;
        RECT -43.630 1521.830 2963.250 1524.930 ;
        RECT -43.630 1341.830 2963.250 1344.930 ;
        RECT -43.630 1161.830 2963.250 1164.930 ;
        RECT -43.630 981.830 2963.250 984.930 ;
        RECT -43.630 801.830 2963.250 804.930 ;
        RECT -43.630 621.830 2963.250 624.930 ;
        RECT -43.630 441.830 2963.250 444.930 ;
        RECT -43.630 261.830 2963.250 264.930 ;
        RECT -43.630 81.830 2963.250 84.930 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.830 17.240 3.150 17.300 ;
        RECT 436.610 17.240 436.930 17.300 ;
        RECT 2.830 17.100 436.930 17.240 ;
        RECT 2.830 17.040 3.150 17.100 ;
        RECT 436.610 17.040 436.930 17.100 ;
      LAYER via ;
        RECT 2.860 17.040 3.120 17.300 ;
        RECT 436.640 17.040 436.900 17.300 ;
      LAYER met2 ;
        RECT 436.430 500.000 436.710 504.000 ;
        RECT 436.470 498.680 436.610 500.000 ;
        RECT 436.470 498.540 436.840 498.680 ;
        RECT 436.700 17.330 436.840 498.540 ;
        RECT 2.860 17.010 3.120 17.330 ;
        RECT 436.640 17.010 436.900 17.330 ;
        RECT 2.920 2.400 3.060 17.010 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 435.690 499.700 436.010 499.760 ;
        RECT 436.840 499.700 437.160 499.760 ;
        RECT 435.690 499.560 437.160 499.700 ;
        RECT 435.690 499.500 436.010 499.560 ;
        RECT 436.840 499.500 437.160 499.560 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 435.690 17.580 436.010 17.640 ;
        RECT 8.350 17.440 436.010 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 435.690 17.380 436.010 17.440 ;
      LAYER via ;
        RECT 435.720 499.500 435.980 499.760 ;
        RECT 436.870 499.500 437.130 499.760 ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 435.720 17.380 435.980 17.640 ;
      LAYER met2 ;
        RECT 436.890 500.000 437.170 504.000 ;
        RECT 436.930 499.790 437.070 500.000 ;
        RECT 435.720 499.470 435.980 499.790 ;
        RECT 436.870 499.470 437.130 499.790 ;
        RECT 435.780 17.670 435.920 499.470 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 435.720 17.350 435.980 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 436.150 491.540 436.470 491.600 ;
        RECT 437.070 491.540 437.390 491.600 ;
        RECT 436.150 491.400 437.390 491.540 ;
        RECT 436.150 491.340 436.470 491.400 ;
        RECT 437.070 491.340 437.390 491.400 ;
        RECT 14.330 17.920 14.650 17.980 ;
        RECT 436.150 17.920 436.470 17.980 ;
        RECT 14.330 17.780 436.470 17.920 ;
        RECT 14.330 17.720 14.650 17.780 ;
        RECT 436.150 17.720 436.470 17.780 ;
      LAYER via ;
        RECT 436.180 491.340 436.440 491.600 ;
        RECT 437.100 491.340 437.360 491.600 ;
        RECT 14.360 17.720 14.620 17.980 ;
        RECT 436.180 17.720 436.440 17.980 ;
      LAYER met2 ;
        RECT 437.350 500.000 437.630 504.000 ;
        RECT 437.390 499.020 437.530 500.000 ;
        RECT 437.160 498.880 437.530 499.020 ;
        RECT 437.160 491.630 437.300 498.880 ;
        RECT 436.180 491.310 436.440 491.630 ;
        RECT 437.100 491.310 437.360 491.630 ;
        RECT 436.240 18.010 436.380 491.310 ;
        RECT 14.360 17.690 14.620 18.010 ;
        RECT 436.180 17.690 436.440 18.010 ;
        RECT 14.420 2.400 14.560 17.690 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 38.250 18.600 38.570 18.660 ;
        RECT 439.830 18.600 440.150 18.660 ;
        RECT 38.250 18.460 440.150 18.600 ;
        RECT 38.250 18.400 38.570 18.460 ;
        RECT 439.830 18.400 440.150 18.460 ;
      LAYER via ;
        RECT 38.280 18.400 38.540 18.660 ;
        RECT 439.860 18.400 440.120 18.660 ;
      LAYER met2 ;
        RECT 439.190 500.000 439.470 504.000 ;
        RECT 439.230 498.850 439.370 500.000 ;
        RECT 439.230 498.710 439.600 498.850 ;
        RECT 439.460 487.970 439.600 498.710 ;
        RECT 439.460 487.830 440.060 487.970 ;
        RECT 439.920 18.690 440.060 487.830 ;
        RECT 38.280 18.370 38.540 18.690 ;
        RECT 439.860 18.370 440.120 18.690 ;
        RECT 38.340 2.400 38.480 18.370 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 453.630 489.840 453.950 489.900 ;
        RECT 454.550 489.840 454.870 489.900 ;
        RECT 453.630 489.700 454.870 489.840 ;
        RECT 453.630 489.640 453.950 489.700 ;
        RECT 454.550 489.640 454.870 489.700 ;
        RECT 239.270 19.280 239.590 19.340 ;
        RECT 452.710 19.280 453.030 19.340 ;
        RECT 239.270 19.140 453.030 19.280 ;
        RECT 239.270 19.080 239.590 19.140 ;
        RECT 452.710 19.080 453.030 19.140 ;
      LAYER via ;
        RECT 453.660 489.640 453.920 489.900 ;
        RECT 454.580 489.640 454.840 489.900 ;
        RECT 239.300 19.080 239.560 19.340 ;
        RECT 452.740 19.080 453.000 19.340 ;
      LAYER met2 ;
        RECT 454.830 500.000 455.110 504.000 ;
        RECT 454.870 498.680 455.010 500.000 ;
        RECT 454.640 498.540 455.010 498.680 ;
        RECT 454.640 489.930 454.780 498.540 ;
        RECT 453.660 489.610 453.920 489.930 ;
        RECT 454.580 489.610 454.840 489.930 ;
        RECT 453.720 473.010 453.860 489.610 ;
        RECT 452.800 472.870 453.860 473.010 ;
        RECT 452.800 19.370 452.940 472.870 ;
        RECT 239.300 19.050 239.560 19.370 ;
        RECT 452.740 19.050 453.000 19.370 ;
        RECT 239.360 2.400 239.500 19.050 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.160 499.160 456.480 499.420 ;
        RECT 456.250 498.400 456.390 499.160 ;
        RECT 455.930 498.200 456.390 498.400 ;
        RECT 455.930 498.140 456.250 498.200 ;
        RECT 455.930 488.820 456.250 488.880 ;
        RECT 459.610 488.820 459.930 488.880 ;
        RECT 455.930 488.680 459.930 488.820 ;
        RECT 455.930 488.620 456.250 488.680 ;
        RECT 459.610 488.620 459.930 488.680 ;
        RECT 256.750 19.960 257.070 20.020 ;
        RECT 460.070 19.960 460.390 20.020 ;
        RECT 256.750 19.820 460.390 19.960 ;
        RECT 256.750 19.760 257.070 19.820 ;
        RECT 460.070 19.760 460.390 19.820 ;
      LAYER via ;
        RECT 456.190 499.160 456.450 499.420 ;
        RECT 455.960 498.140 456.220 498.400 ;
        RECT 455.960 488.620 456.220 488.880 ;
        RECT 459.640 488.620 459.900 488.880 ;
        RECT 256.780 19.760 257.040 20.020 ;
        RECT 460.100 19.760 460.360 20.020 ;
      LAYER met2 ;
        RECT 456.210 500.000 456.490 504.000 ;
        RECT 456.250 499.450 456.390 500.000 ;
        RECT 456.190 499.130 456.450 499.450 ;
        RECT 455.960 498.110 456.220 498.430 ;
        RECT 456.020 488.910 456.160 498.110 ;
        RECT 455.960 488.590 456.220 488.910 ;
        RECT 459.640 488.590 459.900 488.910 ;
        RECT 459.700 473.010 459.840 488.590 ;
        RECT 459.700 472.870 460.300 473.010 ;
        RECT 460.160 20.050 460.300 472.870 ;
        RECT 256.780 19.730 257.040 20.050 ;
        RECT 460.100 19.730 460.360 20.050 ;
        RECT 256.840 2.400 256.980 19.730 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.390 487.460 456.710 487.520 ;
        RECT 457.770 487.460 458.090 487.520 ;
        RECT 456.390 487.320 458.090 487.460 ;
        RECT 456.390 487.260 456.710 487.320 ;
        RECT 457.770 487.260 458.090 487.320 ;
        RECT 274.690 20.300 275.010 20.360 ;
        RECT 456.390 20.300 456.710 20.360 ;
        RECT 274.690 20.160 456.710 20.300 ;
        RECT 274.690 20.100 275.010 20.160 ;
        RECT 456.390 20.100 456.710 20.160 ;
      LAYER via ;
        RECT 456.420 487.260 456.680 487.520 ;
        RECT 457.800 487.260 458.060 487.520 ;
        RECT 274.720 20.100 274.980 20.360 ;
        RECT 456.420 20.100 456.680 20.360 ;
      LAYER met2 ;
        RECT 457.590 500.000 457.870 504.000 ;
        RECT 457.630 499.360 457.770 500.000 ;
        RECT 457.400 499.220 457.770 499.360 ;
        RECT 457.400 498.850 457.540 499.220 ;
        RECT 457.400 498.710 457.770 498.850 ;
        RECT 457.630 498.680 457.770 498.710 ;
        RECT 457.630 498.540 458.000 498.680 ;
        RECT 457.860 487.550 458.000 498.540 ;
        RECT 456.420 487.230 456.680 487.550 ;
        RECT 457.800 487.230 458.060 487.550 ;
        RECT 456.480 20.390 456.620 487.230 ;
        RECT 274.720 20.070 274.980 20.390 ;
        RECT 456.420 20.070 456.680 20.390 ;
        RECT 274.780 2.400 274.920 20.070 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 458.920 499.360 459.240 499.420 ;
        RECT 458.920 499.220 460.300 499.360 ;
        RECT 458.920 499.160 459.240 499.220 ;
        RECT 460.160 496.980 460.300 499.220 ;
        RECT 460.990 496.980 461.310 497.040 ;
        RECT 460.160 496.840 461.310 496.980 ;
        RECT 460.990 496.780 461.310 496.840 ;
        RECT 292.170 20.640 292.490 20.700 ;
        RECT 460.990 20.640 461.310 20.700 ;
        RECT 292.170 20.500 461.310 20.640 ;
        RECT 292.170 20.440 292.490 20.500 ;
        RECT 460.990 20.440 461.310 20.500 ;
      LAYER via ;
        RECT 458.950 499.160 459.210 499.420 ;
        RECT 461.020 496.780 461.280 497.040 ;
        RECT 292.200 20.440 292.460 20.700 ;
        RECT 461.020 20.440 461.280 20.700 ;
      LAYER met2 ;
        RECT 458.970 500.000 459.250 504.000 ;
        RECT 459.010 499.450 459.150 500.000 ;
        RECT 458.950 499.130 459.210 499.450 ;
        RECT 461.020 496.750 461.280 497.070 ;
        RECT 461.080 20.730 461.220 496.750 ;
        RECT 292.200 20.410 292.460 20.730 ;
        RECT 461.020 20.410 461.280 20.730 ;
        RECT 292.260 2.400 292.400 20.410 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 460.300 499.700 460.620 499.760 ;
        RECT 460.300 499.560 460.990 499.700 ;
        RECT 460.300 499.500 460.620 499.560 ;
        RECT 460.850 498.000 460.990 499.560 ;
        RECT 461.450 498.000 461.770 498.060 ;
        RECT 460.850 497.860 461.770 498.000 ;
        RECT 461.450 497.800 461.770 497.860 ;
        RECT 456.850 471.820 457.170 471.880 ;
        RECT 461.450 471.820 461.770 471.880 ;
        RECT 456.850 471.680 461.770 471.820 ;
        RECT 456.850 471.620 457.170 471.680 ;
        RECT 461.450 471.620 461.770 471.680 ;
        RECT 310.110 16.900 310.430 16.960 ;
        RECT 456.850 16.900 457.170 16.960 ;
        RECT 310.110 16.760 457.170 16.900 ;
        RECT 310.110 16.700 310.430 16.760 ;
        RECT 456.850 16.700 457.170 16.760 ;
      LAYER via ;
        RECT 460.330 499.500 460.590 499.760 ;
        RECT 461.480 497.800 461.740 498.060 ;
        RECT 456.880 471.620 457.140 471.880 ;
        RECT 461.480 471.620 461.740 471.880 ;
        RECT 310.140 16.700 310.400 16.960 ;
        RECT 456.880 16.700 457.140 16.960 ;
      LAYER met2 ;
        RECT 460.350 500.000 460.630 504.000 ;
        RECT 460.390 499.790 460.530 500.000 ;
        RECT 460.330 499.470 460.590 499.790 ;
        RECT 461.480 497.770 461.740 498.090 ;
        RECT 461.540 471.910 461.680 497.770 ;
        RECT 456.880 471.590 457.140 471.910 ;
        RECT 461.480 471.590 461.740 471.910 ;
        RECT 456.940 16.990 457.080 471.590 ;
        RECT 310.140 16.670 310.400 16.990 ;
        RECT 456.880 16.670 457.140 16.990 ;
        RECT 310.200 2.400 310.340 16.670 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 461.680 499.500 462.000 499.760 ;
        RECT 461.770 499.360 461.910 499.500 ;
        RECT 461.540 499.220 461.910 499.360 ;
        RECT 461.540 498.340 461.680 499.220 ;
        RECT 461.910 498.340 462.230 498.400 ;
        RECT 461.540 498.200 462.230 498.340 ;
        RECT 461.910 498.140 462.230 498.200 ;
        RECT 457.310 472.160 457.630 472.220 ;
        RECT 461.910 472.160 462.230 472.220 ;
        RECT 457.310 472.020 462.230 472.160 ;
        RECT 457.310 471.960 457.630 472.020 ;
        RECT 461.910 471.960 462.230 472.020 ;
        RECT 327.590 16.560 327.910 16.620 ;
        RECT 457.310 16.560 457.630 16.620 ;
        RECT 327.590 16.420 457.630 16.560 ;
        RECT 327.590 16.360 327.910 16.420 ;
        RECT 457.310 16.360 457.630 16.420 ;
      LAYER via ;
        RECT 461.710 499.500 461.970 499.760 ;
        RECT 461.940 498.140 462.200 498.400 ;
        RECT 457.340 471.960 457.600 472.220 ;
        RECT 461.940 471.960 462.200 472.220 ;
        RECT 327.620 16.360 327.880 16.620 ;
        RECT 457.340 16.360 457.600 16.620 ;
      LAYER met2 ;
        RECT 461.730 500.000 462.010 504.000 ;
        RECT 461.770 499.790 461.910 500.000 ;
        RECT 461.710 499.470 461.970 499.790 ;
        RECT 461.940 498.110 462.200 498.430 ;
        RECT 462.000 472.250 462.140 498.110 ;
        RECT 457.340 471.930 457.600 472.250 ;
        RECT 461.940 471.930 462.200 472.250 ;
        RECT 457.400 16.650 457.540 471.930 ;
        RECT 327.620 16.330 327.880 16.650 ;
        RECT 457.340 16.330 457.600 16.650 ;
        RECT 327.680 2.400 327.820 16.330 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 345.530 16.220 345.850 16.280 ;
        RECT 466.970 16.220 467.290 16.280 ;
        RECT 345.530 16.080 467.290 16.220 ;
        RECT 345.530 16.020 345.850 16.080 ;
        RECT 466.970 16.020 467.290 16.080 ;
      LAYER via ;
        RECT 345.560 16.020 345.820 16.280 ;
        RECT 467.000 16.020 467.260 16.280 ;
      LAYER met2 ;
        RECT 463.110 500.000 463.390 504.000 ;
        RECT 463.150 499.645 463.290 500.000 ;
        RECT 463.080 499.275 463.360 499.645 ;
        RECT 466.990 497.915 467.270 498.285 ;
        RECT 467.060 16.310 467.200 497.915 ;
        RECT 345.560 15.990 345.820 16.310 ;
        RECT 467.000 15.990 467.260 16.310 ;
        RECT 345.620 2.400 345.760 15.990 ;
        RECT 345.410 -4.800 345.970 2.400 ;
      LAYER via2 ;
        RECT 463.080 499.320 463.360 499.600 ;
        RECT 466.990 497.960 467.270 498.240 ;
      LAYER met3 ;
        RECT 463.055 499.610 463.385 499.625 ;
        RECT 461.230 499.310 463.385 499.610 ;
        RECT 461.230 498.250 461.530 499.310 ;
        RECT 463.055 499.295 463.385 499.310 ;
        RECT 466.965 498.250 467.295 498.265 ;
        RECT 461.230 497.950 467.295 498.250 ;
        RECT 466.965 497.935 467.295 497.950 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 358.870 487.800 359.190 487.860 ;
        RECT 464.210 487.800 464.530 487.860 ;
        RECT 358.870 487.660 464.530 487.800 ;
        RECT 358.870 487.600 359.190 487.660 ;
        RECT 464.210 487.600 464.530 487.660 ;
      LAYER via ;
        RECT 358.900 487.600 359.160 487.860 ;
        RECT 464.240 487.600 464.500 487.860 ;
      LAYER met2 ;
        RECT 464.490 500.000 464.770 504.000 ;
        RECT 464.530 499.360 464.670 500.000 ;
        RECT 464.530 499.220 464.900 499.360 ;
        RECT 464.760 497.490 464.900 499.220 ;
        RECT 464.300 497.350 464.900 497.490 ;
        RECT 464.300 487.890 464.440 497.350 ;
        RECT 358.900 487.570 359.160 487.890 ;
        RECT 464.240 487.570 464.500 487.890 ;
        RECT 358.960 82.870 359.100 487.570 ;
        RECT 358.960 82.730 363.240 82.870 ;
        RECT 363.100 2.400 363.240 82.730 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 379.570 479.980 379.890 480.040 ;
        RECT 466.050 479.980 466.370 480.040 ;
        RECT 379.570 479.840 466.370 479.980 ;
        RECT 379.570 479.780 379.890 479.840 ;
        RECT 466.050 479.780 466.370 479.840 ;
      LAYER via ;
        RECT 379.600 479.780 379.860 480.040 ;
        RECT 466.080 479.780 466.340 480.040 ;
      LAYER met2 ;
        RECT 465.870 500.000 466.150 504.000 ;
        RECT 465.910 499.700 466.050 500.000 ;
        RECT 465.680 499.560 466.050 499.700 ;
        RECT 465.680 488.480 465.820 499.560 ;
        RECT 465.680 488.340 466.280 488.480 ;
        RECT 466.140 480.070 466.280 488.340 ;
        RECT 379.600 479.750 379.860 480.070 ;
        RECT 466.080 479.750 466.340 480.070 ;
        RECT 379.660 1.770 379.800 479.750 ;
        RECT 380.830 1.770 381.390 2.400 ;
        RECT 379.660 1.630 381.390 1.770 ;
        RECT 380.830 -4.800 381.390 1.630 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 398.430 30.160 398.750 30.220 ;
        RECT 467.890 30.160 468.210 30.220 ;
        RECT 398.430 30.020 468.210 30.160 ;
        RECT 398.430 29.960 398.750 30.020 ;
        RECT 467.890 29.960 468.210 30.020 ;
      LAYER via ;
        RECT 398.460 29.960 398.720 30.220 ;
        RECT 467.920 29.960 468.180 30.220 ;
      LAYER met2 ;
        RECT 467.250 500.000 467.530 504.000 ;
        RECT 467.290 499.815 467.430 500.000 ;
        RECT 467.220 499.445 467.500 499.815 ;
        RECT 467.450 498.850 467.730 498.965 ;
        RECT 467.450 498.710 468.120 498.850 ;
        RECT 467.450 498.595 467.730 498.710 ;
        RECT 467.980 30.250 468.120 498.710 ;
        RECT 398.460 29.930 398.720 30.250 ;
        RECT 467.920 29.930 468.180 30.250 ;
        RECT 398.520 2.400 398.660 29.930 ;
        RECT 398.310 -4.800 398.870 2.400 ;
      LAYER via2 ;
        RECT 467.220 499.490 467.500 499.770 ;
        RECT 467.450 498.640 467.730 498.920 ;
      LAYER met3 ;
        RECT 467.195 499.465 467.525 499.795 ;
        RECT 467.210 498.945 467.510 499.465 ;
        RECT 467.210 498.630 467.755 498.945 ;
        RECT 467.425 498.615 467.755 498.630 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 55.270 486.440 55.590 486.500 ;
        RECT 440.750 486.440 441.070 486.500 ;
        RECT 55.270 486.300 441.070 486.440 ;
        RECT 55.270 486.240 55.590 486.300 ;
        RECT 440.750 486.240 441.070 486.300 ;
        RECT 55.270 16.900 55.590 16.960 ;
        RECT 59.870 16.900 60.190 16.960 ;
        RECT 55.270 16.760 60.190 16.900 ;
        RECT 55.270 16.700 55.590 16.760 ;
        RECT 59.870 16.700 60.190 16.760 ;
      LAYER via ;
        RECT 55.300 486.240 55.560 486.500 ;
        RECT 440.780 486.240 441.040 486.500 ;
        RECT 55.300 16.700 55.560 16.960 ;
        RECT 59.900 16.700 60.160 16.960 ;
      LAYER met2 ;
        RECT 441.030 500.000 441.310 504.000 ;
        RECT 441.070 498.680 441.210 500.000 ;
        RECT 440.840 498.540 441.210 498.680 ;
        RECT 440.840 486.530 440.980 498.540 ;
        RECT 55.300 486.210 55.560 486.530 ;
        RECT 440.780 486.210 441.040 486.530 ;
        RECT 55.360 16.990 55.500 486.210 ;
        RECT 55.300 16.670 55.560 16.990 ;
        RECT 59.900 16.670 60.160 16.990 ;
        RECT 59.960 1.770 60.100 16.670 ;
        RECT 61.590 1.770 62.150 2.400 ;
        RECT 59.960 1.630 62.150 1.770 ;
        RECT 61.590 -4.800 62.150 1.630 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 465.590 472.840 465.910 472.900 ;
        RECT 468.350 472.840 468.670 472.900 ;
        RECT 465.590 472.700 468.670 472.840 ;
        RECT 465.590 472.640 465.910 472.700 ;
        RECT 468.350 472.640 468.670 472.700 ;
        RECT 414.070 107.000 414.390 107.060 ;
        RECT 465.590 107.000 465.910 107.060 ;
        RECT 414.070 106.860 465.910 107.000 ;
        RECT 414.070 106.800 414.390 106.860 ;
        RECT 465.590 106.800 465.910 106.860 ;
      LAYER via ;
        RECT 465.620 472.640 465.880 472.900 ;
        RECT 468.380 472.640 468.640 472.900 ;
        RECT 414.100 106.800 414.360 107.060 ;
        RECT 465.620 106.800 465.880 107.060 ;
      LAYER met2 ;
        RECT 468.630 500.000 468.910 504.000 ;
        RECT 468.670 499.645 468.810 500.000 ;
        RECT 468.600 499.275 468.880 499.645 ;
        RECT 468.370 498.595 468.650 498.965 ;
        RECT 468.440 472.930 468.580 498.595 ;
        RECT 465.620 472.610 465.880 472.930 ;
        RECT 468.380 472.610 468.640 472.930 ;
        RECT 465.680 107.090 465.820 472.610 ;
        RECT 414.100 106.770 414.360 107.090 ;
        RECT 465.620 106.770 465.880 107.090 ;
        RECT 414.160 82.870 414.300 106.770 ;
        RECT 414.160 82.730 416.600 82.870 ;
        RECT 416.460 2.400 416.600 82.730 ;
        RECT 416.250 -4.800 416.810 2.400 ;
      LAYER via2 ;
        RECT 468.600 499.320 468.880 499.600 ;
        RECT 468.370 498.640 468.650 498.920 ;
      LAYER met3 ;
        RECT 468.575 499.295 468.905 499.625 ;
        RECT 468.590 498.945 468.890 499.295 ;
        RECT 468.345 498.630 468.890 498.945 ;
        RECT 468.345 498.615 468.675 498.630 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.960 499.500 470.280 499.760 ;
        RECT 470.050 499.080 470.190 499.500 ;
        RECT 469.730 498.880 470.190 499.080 ;
        RECT 469.730 498.820 470.050 498.880 ;
        RECT 427.870 489.160 428.190 489.220 ;
        RECT 469.730 489.160 470.050 489.220 ;
        RECT 427.870 489.020 470.050 489.160 ;
        RECT 427.870 488.960 428.190 489.020 ;
        RECT 469.730 488.960 470.050 489.020 ;
      LAYER via ;
        RECT 469.990 499.500 470.250 499.760 ;
        RECT 469.760 498.820 470.020 499.080 ;
        RECT 427.900 488.960 428.160 489.220 ;
        RECT 469.760 488.960 470.020 489.220 ;
      LAYER met2 ;
        RECT 470.010 500.000 470.290 504.000 ;
        RECT 470.050 499.790 470.190 500.000 ;
        RECT 469.990 499.470 470.250 499.790 ;
        RECT 469.760 498.790 470.020 499.110 ;
        RECT 469.820 489.250 469.960 498.790 ;
        RECT 427.900 488.930 428.160 489.250 ;
        RECT 469.760 488.930 470.020 489.250 ;
        RECT 427.960 82.870 428.100 488.930 ;
        RECT 427.960 82.730 430.860 82.870 ;
        RECT 430.720 2.450 430.860 82.730 ;
        RECT 430.720 2.310 432.240 2.450 ;
        RECT 432.100 1.770 432.240 2.310 ;
        RECT 434.190 1.770 434.750 2.400 ;
        RECT 432.100 1.630 434.750 1.770 ;
        RECT 434.190 -4.800 434.750 1.630 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 471.340 498.820 471.660 499.080 ;
        RECT 471.430 498.060 471.570 498.820 ;
        RECT 471.110 497.860 471.570 498.060 ;
        RECT 471.110 497.800 471.430 497.860 ;
        RECT 466.510 484.740 466.830 484.800 ;
        RECT 471.110 484.740 471.430 484.800 ;
        RECT 466.510 484.600 471.430 484.740 ;
        RECT 466.510 484.540 466.830 484.600 ;
        RECT 471.110 484.540 471.430 484.600 ;
        RECT 451.790 15.540 452.110 15.600 ;
        RECT 466.050 15.540 466.370 15.600 ;
        RECT 451.790 15.400 466.370 15.540 ;
        RECT 451.790 15.340 452.110 15.400 ;
        RECT 466.050 15.340 466.370 15.400 ;
      LAYER via ;
        RECT 471.370 498.820 471.630 499.080 ;
        RECT 471.140 497.800 471.400 498.060 ;
        RECT 466.540 484.540 466.800 484.800 ;
        RECT 471.140 484.540 471.400 484.800 ;
        RECT 451.820 15.340 452.080 15.600 ;
        RECT 466.080 15.340 466.340 15.600 ;
      LAYER met2 ;
        RECT 471.390 500.000 471.670 504.000 ;
        RECT 471.430 499.110 471.570 500.000 ;
        RECT 471.370 498.790 471.630 499.110 ;
        RECT 471.140 497.770 471.400 498.090 ;
        RECT 471.200 484.830 471.340 497.770 ;
        RECT 466.540 484.510 466.800 484.830 ;
        RECT 471.140 484.510 471.400 484.830 ;
        RECT 466.600 448.570 466.740 484.510 ;
        RECT 466.140 448.430 466.740 448.570 ;
        RECT 466.140 15.630 466.280 448.430 ;
        RECT 451.820 15.310 452.080 15.630 ;
        RECT 466.080 15.310 466.340 15.630 ;
        RECT 451.880 2.400 452.020 15.310 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 472.720 499.500 473.040 499.760 ;
        RECT 472.810 499.020 472.950 499.500 ;
        RECT 472.810 498.880 473.180 499.020 ;
        RECT 473.040 498.060 473.180 498.880 ;
        RECT 472.950 497.800 473.270 498.060 ;
        RECT 472.950 488.140 473.270 488.200 ;
        RECT 474.330 488.140 474.650 488.200 ;
        RECT 472.950 488.000 474.650 488.140 ;
        RECT 472.950 487.940 473.270 488.000 ;
        RECT 474.330 487.940 474.650 488.000 ;
        RECT 471.570 17.580 471.890 17.640 ;
        RECT 474.330 17.580 474.650 17.640 ;
        RECT 471.570 17.440 474.650 17.580 ;
        RECT 471.570 17.380 471.890 17.440 ;
        RECT 474.330 17.380 474.650 17.440 ;
      LAYER via ;
        RECT 472.750 499.500 473.010 499.760 ;
        RECT 472.980 497.800 473.240 498.060 ;
        RECT 472.980 487.940 473.240 488.200 ;
        RECT 474.360 487.940 474.620 488.200 ;
        RECT 471.600 17.380 471.860 17.640 ;
        RECT 474.360 17.380 474.620 17.640 ;
      LAYER met2 ;
        RECT 472.770 500.000 473.050 504.000 ;
        RECT 472.810 499.790 472.950 500.000 ;
        RECT 472.750 499.470 473.010 499.790 ;
        RECT 472.980 497.770 473.240 498.090 ;
        RECT 473.040 488.230 473.180 497.770 ;
        RECT 472.980 487.910 473.240 488.230 ;
        RECT 474.360 487.910 474.620 488.230 ;
        RECT 474.420 17.670 474.560 487.910 ;
        RECT 471.600 17.350 471.860 17.670 ;
        RECT 474.360 17.350 474.620 17.670 ;
        RECT 469.610 1.770 470.170 2.400 ;
        RECT 471.660 1.770 471.800 17.350 ;
        RECT 469.610 1.630 471.800 1.770 ;
        RECT 469.610 -4.800 470.170 1.630 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 474.100 499.160 474.420 499.420 ;
        RECT 474.190 497.320 474.330 499.160 ;
        RECT 474.790 497.320 475.110 497.380 ;
        RECT 474.190 497.180 475.110 497.320 ;
        RECT 474.790 497.120 475.110 497.180 ;
        RECT 474.790 17.580 475.110 17.640 ;
        RECT 487.210 17.580 487.530 17.640 ;
        RECT 474.790 17.440 487.530 17.580 ;
        RECT 474.790 17.380 475.110 17.440 ;
        RECT 487.210 17.380 487.530 17.440 ;
      LAYER via ;
        RECT 474.130 499.160 474.390 499.420 ;
        RECT 474.820 497.120 475.080 497.380 ;
        RECT 474.820 17.380 475.080 17.640 ;
        RECT 487.240 17.380 487.500 17.640 ;
      LAYER met2 ;
        RECT 474.150 500.000 474.430 504.000 ;
        RECT 474.190 499.450 474.330 500.000 ;
        RECT 474.130 499.130 474.390 499.450 ;
        RECT 474.820 497.090 475.080 497.410 ;
        RECT 474.880 17.670 475.020 497.090 ;
        RECT 474.820 17.350 475.080 17.670 ;
        RECT 487.240 17.350 487.500 17.670 ;
        RECT 487.300 2.400 487.440 17.350 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 475.480 499.500 475.800 499.760 ;
        RECT 475.570 498.340 475.710 499.500 ;
        RECT 475.570 498.200 475.940 498.340 ;
        RECT 475.800 498.060 475.940 498.200 ;
        RECT 475.710 497.800 476.030 498.060 ;
        RECT 471.570 467.740 471.890 467.800 ;
        RECT 475.710 467.740 476.030 467.800 ;
        RECT 471.570 467.600 476.030 467.740 ;
        RECT 471.570 467.540 471.890 467.600 ;
        RECT 475.710 467.540 476.030 467.600 ;
        RECT 471.570 18.940 471.890 19.000 ;
        RECT 505.150 18.940 505.470 19.000 ;
        RECT 471.570 18.800 505.470 18.940 ;
        RECT 471.570 18.740 471.890 18.800 ;
        RECT 505.150 18.740 505.470 18.800 ;
      LAYER via ;
        RECT 475.510 499.500 475.770 499.760 ;
        RECT 475.740 497.800 476.000 498.060 ;
        RECT 471.600 467.540 471.860 467.800 ;
        RECT 475.740 467.540 476.000 467.800 ;
        RECT 471.600 18.740 471.860 19.000 ;
        RECT 505.180 18.740 505.440 19.000 ;
      LAYER met2 ;
        RECT 475.530 500.000 475.810 504.000 ;
        RECT 475.570 499.790 475.710 500.000 ;
        RECT 475.510 499.470 475.770 499.790 ;
        RECT 475.740 497.770 476.000 498.090 ;
        RECT 475.800 467.830 475.940 497.770 ;
        RECT 471.600 467.510 471.860 467.830 ;
        RECT 475.740 467.510 476.000 467.830 ;
        RECT 471.660 19.030 471.800 467.510 ;
        RECT 471.600 18.710 471.860 19.030 ;
        RECT 505.180 18.710 505.440 19.030 ;
        RECT 505.240 2.400 505.380 18.710 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 477.090 16.560 477.410 16.620 ;
        RECT 522.630 16.560 522.950 16.620 ;
        RECT 477.090 16.420 522.950 16.560 ;
        RECT 477.090 16.360 477.410 16.420 ;
        RECT 522.630 16.360 522.950 16.420 ;
      LAYER via ;
        RECT 477.120 16.360 477.380 16.620 ;
        RECT 522.660 16.360 522.920 16.620 ;
      LAYER met2 ;
        RECT 476.910 500.000 477.190 504.000 ;
        RECT 476.950 499.645 477.090 500.000 ;
        RECT 476.880 499.275 477.160 499.645 ;
        RECT 477.110 498.595 477.390 498.965 ;
        RECT 477.180 16.650 477.320 498.595 ;
        RECT 477.120 16.330 477.380 16.650 ;
        RECT 522.660 16.330 522.920 16.650 ;
        RECT 522.720 2.400 522.860 16.330 ;
        RECT 522.510 -4.800 523.070 2.400 ;
      LAYER via2 ;
        RECT 476.880 499.320 477.160 499.600 ;
        RECT 477.110 498.640 477.390 498.920 ;
      LAYER met3 ;
        RECT 476.855 499.295 477.185 499.625 ;
        RECT 476.870 498.945 477.170 499.295 ;
        RECT 476.870 498.630 477.415 498.945 ;
        RECT 477.085 498.615 477.415 498.630 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 478.240 499.700 478.560 499.760 ;
        RECT 478.240 499.560 479.850 499.700 ;
        RECT 478.240 499.500 478.560 499.560 ;
        RECT 479.710 497.320 479.850 499.560 ;
        RECT 481.690 497.320 482.010 497.380 ;
        RECT 479.710 497.180 482.010 497.320 ;
        RECT 481.690 497.120 482.010 497.180 ;
        RECT 481.690 16.900 482.010 16.960 ;
        RECT 540.570 16.900 540.890 16.960 ;
        RECT 481.690 16.760 540.890 16.900 ;
        RECT 481.690 16.700 482.010 16.760 ;
        RECT 540.570 16.700 540.890 16.760 ;
      LAYER via ;
        RECT 478.270 499.500 478.530 499.760 ;
        RECT 481.720 497.120 481.980 497.380 ;
        RECT 481.720 16.700 481.980 16.960 ;
        RECT 540.600 16.700 540.860 16.960 ;
      LAYER met2 ;
        RECT 478.290 500.000 478.570 504.000 ;
        RECT 478.330 499.790 478.470 500.000 ;
        RECT 478.270 499.470 478.530 499.790 ;
        RECT 481.720 497.090 481.980 497.410 ;
        RECT 481.780 483.070 481.920 497.090 ;
        RECT 481.780 482.930 482.380 483.070 ;
        RECT 482.240 420.970 482.380 482.930 ;
        RECT 481.780 420.830 482.380 420.970 ;
        RECT 481.780 16.990 481.920 420.830 ;
        RECT 481.720 16.670 481.980 16.990 ;
        RECT 540.600 16.670 540.860 16.990 ;
        RECT 540.660 2.400 540.800 16.670 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 479.620 500.180 479.940 500.440 ;
        RECT 479.710 500.040 479.850 500.180 ;
        RECT 477.870 499.900 479.850 500.040 ;
        RECT 477.870 497.720 478.010 499.900 ;
        RECT 477.550 497.520 478.010 497.720 ;
        RECT 477.550 497.460 477.870 497.520 ;
        RECT 477.550 19.280 477.870 19.340 ;
        RECT 499.630 19.280 499.950 19.340 ;
        RECT 477.550 19.140 499.950 19.280 ;
        RECT 477.550 19.080 477.870 19.140 ;
        RECT 499.630 19.080 499.950 19.140 ;
        RECT 499.630 17.920 499.950 17.980 ;
        RECT 558.050 17.920 558.370 17.980 ;
        RECT 499.630 17.780 558.370 17.920 ;
        RECT 499.630 17.720 499.950 17.780 ;
        RECT 558.050 17.720 558.370 17.780 ;
      LAYER via ;
        RECT 479.650 500.180 479.910 500.440 ;
        RECT 477.580 497.460 477.840 497.720 ;
        RECT 477.580 19.080 477.840 19.340 ;
        RECT 499.660 19.080 499.920 19.340 ;
        RECT 499.660 17.720 499.920 17.980 ;
        RECT 558.080 17.720 558.340 17.980 ;
      LAYER met2 ;
        RECT 479.670 500.470 479.950 504.000 ;
        RECT 479.650 500.150 479.950 500.470 ;
        RECT 479.670 500.000 479.950 500.150 ;
        RECT 477.580 497.430 477.840 497.750 ;
        RECT 477.640 19.370 477.780 497.430 ;
        RECT 477.580 19.050 477.840 19.370 ;
        RECT 499.660 19.050 499.920 19.370 ;
        RECT 499.720 18.010 499.860 19.050 ;
        RECT 499.660 17.690 499.920 18.010 ;
        RECT 558.080 17.690 558.340 18.010 ;
        RECT 558.140 2.400 558.280 17.690 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 481.000 499.500 481.320 499.760 ;
        RECT 481.090 499.080 481.230 499.500 ;
        RECT 481.000 498.820 481.320 499.080 ;
      LAYER via ;
        RECT 481.030 499.500 481.290 499.760 ;
        RECT 481.030 498.820 481.290 499.080 ;
      LAYER met2 ;
        RECT 481.050 500.000 481.330 504.000 ;
        RECT 481.090 499.790 481.230 500.000 ;
        RECT 481.030 499.470 481.290 499.790 ;
        RECT 481.030 498.965 481.290 499.110 ;
        RECT 481.020 498.595 481.300 498.965 ;
        RECT 576.010 23.955 576.290 24.325 ;
        RECT 576.080 2.400 576.220 23.955 ;
        RECT 575.870 -4.800 576.430 2.400 ;
      LAYER via2 ;
        RECT 481.020 498.640 481.300 498.920 ;
        RECT 576.010 24.000 576.290 24.280 ;
      LAYER met3 ;
        RECT 478.670 498.930 479.050 498.940 ;
        RECT 480.995 498.930 481.325 498.945 ;
        RECT 478.670 498.630 481.325 498.930 ;
        RECT 478.670 498.620 479.050 498.630 ;
        RECT 480.995 498.615 481.325 498.630 ;
        RECT 478.670 24.290 479.050 24.300 ;
        RECT 575.985 24.290 576.315 24.305 ;
        RECT 478.670 23.990 576.315 24.290 ;
        RECT 478.670 23.980 479.050 23.990 ;
        RECT 575.985 23.975 576.315 23.990 ;
      LAYER via3 ;
        RECT 478.700 498.620 479.020 498.940 ;
        RECT 478.700 23.980 479.020 24.300 ;
      LAYER met4 ;
        RECT 478.695 498.615 479.025 498.945 ;
        RECT 478.710 24.305 479.010 498.615 ;
        RECT 478.695 23.975 479.025 24.305 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.820 499.500 443.140 499.760 ;
        RECT 442.910 498.060 443.050 499.500 ;
        RECT 442.590 497.860 443.050 498.060 ;
        RECT 442.590 497.800 442.910 497.860 ;
      LAYER via ;
        RECT 442.850 499.500 443.110 499.760 ;
        RECT 442.620 497.800 442.880 498.060 ;
      LAYER met2 ;
        RECT 442.870 500.000 443.150 504.000 ;
        RECT 442.910 499.790 443.050 500.000 ;
        RECT 442.850 499.470 443.110 499.790 ;
        RECT 442.620 497.770 442.880 498.090 ;
        RECT 442.680 492.845 442.820 497.770 ;
        RECT 442.610 492.475 442.890 492.845 ;
        RECT 85.190 24.635 85.470 25.005 ;
        RECT 85.260 2.400 85.400 24.635 ;
        RECT 85.050 -4.800 85.610 2.400 ;
      LAYER via2 ;
        RECT 442.610 492.520 442.890 492.800 ;
        RECT 85.190 24.680 85.470 24.960 ;
      LAYER met3 ;
        RECT 442.585 492.820 442.915 492.825 ;
        RECT 442.585 492.810 443.170 492.820 ;
        RECT 442.585 492.510 443.370 492.810 ;
        RECT 442.585 492.500 443.170 492.510 ;
        RECT 442.585 492.495 442.915 492.500 ;
        RECT 85.165 24.970 85.495 24.985 ;
        RECT 442.790 24.970 443.170 24.980 ;
        RECT 85.165 24.670 443.170 24.970 ;
        RECT 85.165 24.655 85.495 24.670 ;
        RECT 442.790 24.660 443.170 24.670 ;
      LAYER via3 ;
        RECT 442.820 492.500 443.140 492.820 ;
        RECT 442.820 24.660 443.140 24.980 ;
      LAYER met4 ;
        RECT 442.815 492.495 443.145 492.825 ;
        RECT 442.830 24.985 443.130 492.495 ;
        RECT 442.815 24.655 443.145 24.985 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 482.610 487.120 482.930 487.180 ;
        RECT 556.670 487.120 556.990 487.180 ;
        RECT 482.610 486.980 556.990 487.120 ;
        RECT 482.610 486.920 482.930 486.980 ;
        RECT 556.670 486.920 556.990 486.980 ;
        RECT 558.510 17.920 558.830 17.980 ;
        RECT 593.930 17.920 594.250 17.980 ;
        RECT 558.510 17.780 594.250 17.920 ;
        RECT 558.510 17.720 558.830 17.780 ;
        RECT 593.930 17.720 594.250 17.780 ;
      LAYER via ;
        RECT 482.640 486.920 482.900 487.180 ;
        RECT 556.700 486.920 556.960 487.180 ;
        RECT 558.540 17.720 558.800 17.980 ;
        RECT 593.960 17.720 594.220 17.980 ;
      LAYER met2 ;
        RECT 482.430 500.000 482.710 504.000 ;
        RECT 482.470 498.680 482.610 500.000 ;
        RECT 482.470 498.540 482.840 498.680 ;
        RECT 482.700 487.210 482.840 498.540 ;
        RECT 482.640 486.890 482.900 487.210 ;
        RECT 556.700 486.890 556.960 487.210 ;
        RECT 556.760 82.870 556.900 486.890 ;
        RECT 556.760 82.730 558.740 82.870 ;
        RECT 558.600 18.010 558.740 82.730 ;
        RECT 558.540 17.690 558.800 18.010 ;
        RECT 593.960 17.690 594.220 18.010 ;
        RECT 594.020 2.400 594.160 17.690 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.530 472.500 483.850 472.560 ;
        RECT 485.830 472.500 486.150 472.560 ;
        RECT 483.530 472.360 486.150 472.500 ;
        RECT 483.530 472.300 483.850 472.360 ;
        RECT 485.830 472.300 486.150 472.360 ;
        RECT 485.830 25.060 486.150 25.120 ;
        RECT 611.410 25.060 611.730 25.120 ;
        RECT 485.830 24.920 611.730 25.060 ;
        RECT 485.830 24.860 486.150 24.920 ;
        RECT 611.410 24.860 611.730 24.920 ;
      LAYER via ;
        RECT 483.560 472.300 483.820 472.560 ;
        RECT 485.860 472.300 486.120 472.560 ;
        RECT 485.860 24.860 486.120 25.120 ;
        RECT 611.440 24.860 611.700 25.120 ;
      LAYER met2 ;
        RECT 483.810 500.000 484.090 504.000 ;
        RECT 483.850 498.340 483.990 500.000 ;
        RECT 483.620 498.200 483.990 498.340 ;
        RECT 483.620 472.590 483.760 498.200 ;
        RECT 483.560 472.270 483.820 472.590 ;
        RECT 485.860 472.270 486.120 472.590 ;
        RECT 485.920 25.150 486.060 472.270 ;
        RECT 485.860 24.830 486.120 25.150 ;
        RECT 611.440 24.830 611.700 25.150 ;
        RECT 611.500 2.400 611.640 24.830 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 444.660 498.820 444.980 499.080 ;
        RECT 443.510 498.340 443.830 498.400 ;
        RECT 444.750 498.340 444.890 498.820 ;
        RECT 443.510 498.200 444.890 498.340 ;
        RECT 443.510 498.140 443.830 498.200 ;
        RECT 109.090 24.380 109.410 24.440 ;
        RECT 443.050 24.380 443.370 24.440 ;
        RECT 109.090 24.240 443.370 24.380 ;
        RECT 109.090 24.180 109.410 24.240 ;
        RECT 443.050 24.180 443.370 24.240 ;
      LAYER via ;
        RECT 444.690 498.820 444.950 499.080 ;
        RECT 443.540 498.140 443.800 498.400 ;
        RECT 109.120 24.180 109.380 24.440 ;
        RECT 443.080 24.180 443.340 24.440 ;
      LAYER met2 ;
        RECT 444.710 500.000 444.990 504.000 ;
        RECT 444.750 499.110 444.890 500.000 ;
        RECT 444.690 498.790 444.950 499.110 ;
        RECT 443.540 498.110 443.800 498.430 ;
        RECT 443.600 491.880 443.740 498.110 ;
        RECT 443.140 491.740 443.740 491.880 ;
        RECT 443.140 24.470 443.280 491.740 ;
        RECT 109.120 24.150 109.380 24.470 ;
        RECT 443.080 24.150 443.340 24.470 ;
        RECT 109.180 2.400 109.320 24.150 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 132.550 25.060 132.870 25.120 ;
        RECT 446.270 25.060 446.590 25.120 ;
        RECT 132.550 24.920 446.590 25.060 ;
        RECT 132.550 24.860 132.870 24.920 ;
        RECT 446.270 24.860 446.590 24.920 ;
      LAYER via ;
        RECT 132.580 24.860 132.840 25.120 ;
        RECT 446.300 24.860 446.560 25.120 ;
      LAYER met2 ;
        RECT 446.550 500.000 446.830 504.000 ;
        RECT 446.590 499.645 446.730 500.000 ;
        RECT 446.520 499.275 446.800 499.645 ;
        RECT 446.290 497.915 446.570 498.285 ;
        RECT 446.360 25.150 446.500 497.915 ;
        RECT 132.580 24.830 132.840 25.150 ;
        RECT 446.300 24.830 446.560 25.150 ;
        RECT 132.640 2.400 132.780 24.830 ;
        RECT 132.430 -4.800 132.990 2.400 ;
      LAYER via2 ;
        RECT 446.520 499.320 446.800 499.600 ;
        RECT 446.290 497.960 446.570 498.240 ;
      LAYER met3 ;
        RECT 446.495 499.295 446.825 499.625 ;
        RECT 446.510 498.265 446.810 499.295 ;
        RECT 446.265 497.950 446.810 498.265 ;
        RECT 446.265 497.935 446.595 497.950 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 447.880 499.500 448.200 499.760 ;
        RECT 447.970 499.080 448.110 499.500 ;
        RECT 447.880 498.820 448.200 499.080 ;
        RECT 443.510 483.040 443.830 483.100 ;
        RECT 448.110 483.040 448.430 483.100 ;
        RECT 443.510 482.900 448.430 483.040 ;
        RECT 443.510 482.840 443.830 482.900 ;
        RECT 448.110 482.840 448.430 482.900 ;
        RECT 150.490 25.400 150.810 25.460 ;
        RECT 443.510 25.400 443.830 25.460 ;
        RECT 150.490 25.260 443.830 25.400 ;
        RECT 150.490 25.200 150.810 25.260 ;
        RECT 443.510 25.200 443.830 25.260 ;
      LAYER via ;
        RECT 447.910 499.500 448.170 499.760 ;
        RECT 447.910 498.820 448.170 499.080 ;
        RECT 443.540 482.840 443.800 483.100 ;
        RECT 448.140 482.840 448.400 483.100 ;
        RECT 150.520 25.200 150.780 25.460 ;
        RECT 443.540 25.200 443.800 25.460 ;
      LAYER met2 ;
        RECT 447.930 500.000 448.210 504.000 ;
        RECT 447.970 499.790 448.110 500.000 ;
        RECT 447.910 499.470 448.170 499.790 ;
        RECT 447.910 498.850 448.170 499.110 ;
        RECT 447.910 498.790 448.340 498.850 ;
        RECT 447.970 498.710 448.340 498.790 ;
        RECT 448.200 483.130 448.340 498.710 ;
        RECT 443.540 482.810 443.800 483.130 ;
        RECT 448.140 482.810 448.400 483.130 ;
        RECT 443.600 25.490 443.740 482.810 ;
        RECT 150.520 25.170 150.780 25.490 ;
        RECT 443.540 25.170 443.800 25.490 ;
        RECT 150.580 2.400 150.720 25.170 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.310 500.000 449.590 504.000 ;
        RECT 449.350 499.815 449.490 500.000 ;
        RECT 449.280 499.445 449.560 499.815 ;
        RECT 167.990 25.315 168.270 25.685 ;
        RECT 168.060 2.400 168.200 25.315 ;
        RECT 167.850 -4.800 168.410 2.400 ;
      LAYER via2 ;
        RECT 449.280 499.490 449.560 499.770 ;
        RECT 167.990 25.360 168.270 25.640 ;
      LAYER met3 ;
        RECT 449.255 499.620 449.585 499.795 ;
        RECT 449.230 499.610 449.610 499.620 ;
        RECT 449.230 499.310 449.870 499.610 ;
        RECT 449.230 499.300 449.610 499.310 ;
        RECT 448.310 449.290 448.690 449.300 ;
        RECT 450.150 449.290 450.530 449.300 ;
        RECT 448.310 448.990 450.530 449.290 ;
        RECT 448.310 448.980 448.690 448.990 ;
        RECT 450.150 448.980 450.530 448.990 ;
        RECT 167.965 25.650 168.295 25.665 ;
        RECT 448.310 25.650 448.690 25.660 ;
        RECT 167.965 25.350 448.690 25.650 ;
        RECT 167.965 25.335 168.295 25.350 ;
        RECT 448.310 25.340 448.690 25.350 ;
      LAYER via3 ;
        RECT 449.260 499.300 449.580 499.620 ;
        RECT 448.340 448.980 448.660 449.300 ;
        RECT 450.180 448.980 450.500 449.300 ;
        RECT 448.340 25.340 448.660 25.660 ;
      LAYER met4 ;
        RECT 449.255 499.610 449.585 499.625 ;
        RECT 449.255 499.310 450.490 499.610 ;
        RECT 449.255 499.295 449.585 499.310 ;
        RECT 450.190 449.305 450.490 499.310 ;
        RECT 448.335 448.975 448.665 449.305 ;
        RECT 450.175 448.975 450.505 449.305 ;
        RECT 448.350 25.665 448.650 448.975 ;
        RECT 448.335 25.335 448.665 25.665 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 185.910 25.740 186.230 25.800 ;
        RECT 450.410 25.740 450.730 25.800 ;
        RECT 185.910 25.600 450.730 25.740 ;
        RECT 185.910 25.540 186.230 25.600 ;
        RECT 450.410 25.540 450.730 25.600 ;
      LAYER via ;
        RECT 185.940 25.540 186.200 25.800 ;
        RECT 450.440 25.540 450.700 25.800 ;
      LAYER met2 ;
        RECT 450.690 500.000 450.970 504.000 ;
        RECT 450.730 499.815 450.870 500.000 ;
        RECT 450.660 499.445 450.940 499.815 ;
        RECT 450.430 498.595 450.710 498.965 ;
        RECT 450.500 25.830 450.640 498.595 ;
        RECT 185.940 25.510 186.200 25.830 ;
        RECT 450.440 25.510 450.700 25.830 ;
        RECT 186.000 2.400 186.140 25.510 ;
        RECT 185.790 -4.800 186.350 2.400 ;
      LAYER via2 ;
        RECT 450.660 499.490 450.940 499.770 ;
        RECT 450.430 498.640 450.710 498.920 ;
      LAYER met3 ;
        RECT 450.635 499.780 450.965 499.795 ;
        RECT 450.635 499.480 451.640 499.780 ;
        RECT 450.635 499.465 450.965 499.480 ;
        RECT 450.405 498.930 450.735 498.945 ;
        RECT 451.340 498.930 451.640 499.480 ;
        RECT 450.405 498.630 451.640 498.930 ;
        RECT 450.405 498.615 450.735 498.630 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 203.390 26.420 203.710 26.480 ;
        RECT 450.870 26.420 451.190 26.480 ;
        RECT 203.390 26.280 451.190 26.420 ;
        RECT 203.390 26.220 203.710 26.280 ;
        RECT 450.870 26.220 451.190 26.280 ;
      LAYER via ;
        RECT 203.420 26.220 203.680 26.480 ;
        RECT 450.900 26.220 451.160 26.480 ;
      LAYER met2 ;
        RECT 452.070 500.000 452.350 504.000 ;
        RECT 452.110 498.170 452.250 500.000 ;
        RECT 451.880 498.030 452.250 498.170 ;
        RECT 451.880 488.140 452.020 498.030 ;
        RECT 451.420 488.000 452.020 488.140 ;
        RECT 451.420 473.010 451.560 488.000 ;
        RECT 450.960 472.870 451.560 473.010 ;
        RECT 450.960 26.510 451.100 472.870 ;
        RECT 203.420 26.190 203.680 26.510 ;
        RECT 450.900 26.190 451.160 26.510 ;
        RECT 203.480 2.400 203.620 26.190 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 453.400 499.500 453.720 499.760 ;
        RECT 449.950 497.320 450.270 497.380 ;
        RECT 453.490 497.320 453.630 499.500 ;
        RECT 449.950 497.180 453.630 497.320 ;
        RECT 449.950 497.120 450.270 497.180 ;
        RECT 221.330 26.760 221.650 26.820 ;
        RECT 449.950 26.760 450.270 26.820 ;
        RECT 221.330 26.620 450.270 26.760 ;
        RECT 221.330 26.560 221.650 26.620 ;
        RECT 449.950 26.560 450.270 26.620 ;
      LAYER via ;
        RECT 453.430 499.500 453.690 499.760 ;
        RECT 449.980 497.120 450.240 497.380 ;
        RECT 221.360 26.560 221.620 26.820 ;
        RECT 449.980 26.560 450.240 26.820 ;
      LAYER met2 ;
        RECT 453.450 500.000 453.730 504.000 ;
        RECT 453.490 499.790 453.630 500.000 ;
        RECT 453.430 499.470 453.690 499.790 ;
        RECT 449.980 497.090 450.240 497.410 ;
        RECT 450.040 26.850 450.180 497.090 ;
        RECT 221.360 26.530 221.620 26.850 ;
        RECT 449.980 26.530 450.240 26.850 ;
        RECT 221.420 2.400 221.560 26.530 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 24.040 20.630 24.100 ;
        RECT 437.530 24.040 437.850 24.100 ;
        RECT 20.310 23.900 437.850 24.040 ;
        RECT 20.310 23.840 20.630 23.900 ;
        RECT 437.530 23.840 437.850 23.900 ;
      LAYER via ;
        RECT 20.340 23.840 20.600 24.100 ;
        RECT 437.560 23.840 437.820 24.100 ;
      LAYER met2 ;
        RECT 437.810 500.000 438.090 504.000 ;
        RECT 437.850 498.680 437.990 500.000 ;
        RECT 437.620 498.540 437.990 498.680 ;
        RECT 437.620 24.130 437.760 498.540 ;
        RECT 20.340 23.810 20.600 24.130 ;
        RECT 437.560 23.810 437.820 24.130 ;
        RECT 20.400 2.400 20.540 23.810 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 43.770 37.980 44.090 38.040 ;
        RECT 437.990 37.980 438.310 38.040 ;
        RECT 43.770 37.840 438.310 37.980 ;
        RECT 43.770 37.780 44.090 37.840 ;
        RECT 437.990 37.780 438.310 37.840 ;
      LAYER via ;
        RECT 43.800 37.780 44.060 38.040 ;
        RECT 438.020 37.780 438.280 38.040 ;
      LAYER met2 ;
        RECT 439.650 500.000 439.930 504.000 ;
        RECT 439.690 499.645 439.830 500.000 ;
        RECT 439.620 499.275 439.900 499.645 ;
        RECT 438.010 491.115 438.290 491.485 ;
        RECT 438.080 38.070 438.220 491.115 ;
        RECT 43.800 37.750 44.060 38.070 ;
        RECT 438.020 37.750 438.280 38.070 ;
        RECT 43.860 2.400 44.000 37.750 ;
        RECT 43.650 -4.800 44.210 2.400 ;
      LAYER via2 ;
        RECT 439.620 499.320 439.900 499.600 ;
        RECT 438.010 491.160 438.290 491.440 ;
      LAYER met3 ;
        RECT 438.190 499.610 438.570 499.620 ;
        RECT 439.595 499.610 439.925 499.625 ;
        RECT 438.190 499.310 439.925 499.610 ;
        RECT 438.190 499.300 438.570 499.310 ;
        RECT 439.595 499.295 439.925 499.310 ;
        RECT 437.985 491.460 438.315 491.465 ;
        RECT 437.985 491.450 438.570 491.460 ;
        RECT 437.760 491.150 438.570 491.450 ;
        RECT 437.985 491.140 438.570 491.150 ;
        RECT 437.985 491.135 438.315 491.140 ;
      LAYER via3 ;
        RECT 438.220 499.300 438.540 499.620 ;
        RECT 438.220 491.140 438.540 491.460 ;
      LAYER met4 ;
        RECT 438.215 499.295 438.545 499.625 ;
        RECT 438.230 491.465 438.530 499.295 ;
        RECT 438.215 491.135 438.545 491.465 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.240 499.500 455.560 499.760 ;
        RECT 455.330 499.360 455.470 499.500 ;
        RECT 455.100 499.220 455.470 499.360 ;
        RECT 455.100 498.060 455.240 499.220 ;
        RECT 455.010 497.800 455.330 498.060 ;
      LAYER via ;
        RECT 455.270 499.500 455.530 499.760 ;
        RECT 455.040 497.800 455.300 498.060 ;
      LAYER met2 ;
        RECT 455.290 500.000 455.570 504.000 ;
        RECT 455.330 499.790 455.470 500.000 ;
        RECT 455.270 499.470 455.530 499.790 ;
        RECT 455.040 497.770 455.300 498.090 ;
        RECT 455.100 489.445 455.240 497.770 ;
        RECT 455.030 489.075 455.310 489.445 ;
        RECT 244.810 30.755 245.090 31.125 ;
        RECT 244.880 2.400 245.020 30.755 ;
        RECT 244.670 -4.800 245.230 2.400 ;
      LAYER via2 ;
        RECT 455.030 489.120 455.310 489.400 ;
        RECT 244.810 30.800 245.090 31.080 ;
      LAYER met3 ;
        RECT 455.005 489.410 455.335 489.425 ;
        RECT 456.590 489.410 456.970 489.420 ;
        RECT 455.005 489.110 456.970 489.410 ;
        RECT 455.005 489.095 455.335 489.110 ;
        RECT 456.590 489.100 456.970 489.110 ;
        RECT 244.785 31.090 245.115 31.105 ;
        RECT 456.590 31.090 456.970 31.100 ;
        RECT 244.785 30.790 456.970 31.090 ;
        RECT 244.785 30.775 245.115 30.790 ;
        RECT 456.590 30.780 456.970 30.790 ;
      LAYER via3 ;
        RECT 456.620 489.100 456.940 489.420 ;
        RECT 456.620 30.780 456.940 31.100 ;
      LAYER met4 ;
        RECT 456.615 489.095 456.945 489.425 ;
        RECT 456.630 31.105 456.930 489.095 ;
        RECT 456.615 30.775 456.945 31.105 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.620 499.020 456.940 499.080 ;
        RECT 456.620 498.820 457.080 499.020 ;
        RECT 456.940 498.060 457.080 498.820 ;
        RECT 456.850 497.800 457.170 498.060 ;
        RECT 262.730 30.840 263.050 30.900 ;
        RECT 457.770 30.840 458.090 30.900 ;
        RECT 262.730 30.700 458.090 30.840 ;
        RECT 262.730 30.640 263.050 30.700 ;
        RECT 457.770 30.640 458.090 30.700 ;
      LAYER via ;
        RECT 456.650 498.820 456.910 499.080 ;
        RECT 456.880 497.800 457.140 498.060 ;
        RECT 262.760 30.640 263.020 30.900 ;
        RECT 457.800 30.640 458.060 30.900 ;
      LAYER met2 ;
        RECT 456.670 500.000 456.950 504.000 ;
        RECT 456.710 499.110 456.850 500.000 ;
        RECT 456.650 498.790 456.910 499.110 ;
        RECT 456.880 497.770 457.140 498.090 ;
        RECT 456.940 473.010 457.080 497.770 ;
        RECT 456.940 472.870 458.000 473.010 ;
        RECT 457.860 30.930 458.000 472.870 ;
        RECT 262.760 30.610 263.020 30.930 ;
        RECT 457.800 30.610 458.060 30.930 ;
        RECT 262.820 2.400 262.960 30.610 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 459.610 472.500 459.930 472.560 ;
        RECT 460.530 472.500 460.850 472.560 ;
        RECT 459.610 472.360 460.850 472.500 ;
        RECT 459.610 472.300 459.930 472.360 ;
        RECT 460.530 472.300 460.850 472.360 ;
        RECT 280.210 31.180 280.530 31.240 ;
        RECT 459.610 31.180 459.930 31.240 ;
        RECT 280.210 31.040 459.930 31.180 ;
        RECT 280.210 30.980 280.530 31.040 ;
        RECT 459.610 30.980 459.930 31.040 ;
      LAYER via ;
        RECT 459.640 472.300 459.900 472.560 ;
        RECT 460.560 472.300 460.820 472.560 ;
        RECT 280.240 30.980 280.500 31.240 ;
        RECT 459.640 30.980 459.900 31.240 ;
      LAYER met2 ;
        RECT 458.050 500.000 458.330 504.000 ;
        RECT 458.090 499.645 458.230 500.000 ;
        RECT 458.020 499.275 458.300 499.645 ;
        RECT 460.090 497.235 460.370 497.605 ;
        RECT 460.160 473.690 460.300 497.235 ;
        RECT 460.160 473.550 460.760 473.690 ;
        RECT 460.620 472.590 460.760 473.550 ;
        RECT 459.640 472.270 459.900 472.590 ;
        RECT 460.560 472.270 460.820 472.590 ;
        RECT 459.700 31.270 459.840 472.270 ;
        RECT 280.240 30.950 280.500 31.270 ;
        RECT 459.640 30.950 459.900 31.270 ;
        RECT 280.300 2.400 280.440 30.950 ;
        RECT 280.090 -4.800 280.650 2.400 ;
      LAYER via2 ;
        RECT 458.020 499.320 458.300 499.600 ;
        RECT 460.090 497.280 460.370 497.560 ;
      LAYER met3 ;
        RECT 457.995 499.610 458.325 499.625 ;
        RECT 457.995 499.310 460.380 499.610 ;
        RECT 457.995 499.295 458.325 499.310 ;
        RECT 460.080 497.585 460.380 499.310 ;
        RECT 460.065 497.255 460.395 497.585 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 459.380 499.700 459.700 499.760 ;
        RECT 458.550 499.560 459.700 499.700 ;
        RECT 458.550 498.000 458.690 499.560 ;
        RECT 459.380 499.500 459.700 499.560 ;
        RECT 459.150 498.000 459.470 498.060 ;
        RECT 458.550 497.860 459.470 498.000 ;
        RECT 459.150 497.800 459.470 497.860 ;
        RECT 298.150 31.860 298.470 31.920 ;
        RECT 459.150 31.860 459.470 31.920 ;
        RECT 298.150 31.720 459.470 31.860 ;
        RECT 298.150 31.660 298.470 31.720 ;
        RECT 459.150 31.660 459.470 31.720 ;
      LAYER via ;
        RECT 459.410 499.500 459.670 499.760 ;
        RECT 459.180 497.800 459.440 498.060 ;
        RECT 298.180 31.660 298.440 31.920 ;
        RECT 459.180 31.660 459.440 31.920 ;
      LAYER met2 ;
        RECT 459.430 500.000 459.710 504.000 ;
        RECT 459.470 499.790 459.610 500.000 ;
        RECT 459.410 499.470 459.670 499.790 ;
        RECT 459.180 497.770 459.440 498.090 ;
        RECT 459.240 31.950 459.380 497.770 ;
        RECT 298.180 31.630 298.440 31.950 ;
        RECT 459.180 31.630 459.440 31.950 ;
        RECT 298.240 2.400 298.380 31.630 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 458.690 474.200 459.010 474.260 ;
        RECT 460.530 474.200 460.850 474.260 ;
        RECT 458.690 474.060 460.850 474.200 ;
        RECT 458.690 474.000 459.010 474.060 ;
        RECT 460.530 474.000 460.850 474.060 ;
        RECT 316.090 32.200 316.410 32.260 ;
        RECT 458.690 32.200 459.010 32.260 ;
        RECT 316.090 32.060 459.010 32.200 ;
        RECT 316.090 32.000 316.410 32.060 ;
        RECT 458.690 32.000 459.010 32.060 ;
      LAYER via ;
        RECT 458.720 474.000 458.980 474.260 ;
        RECT 460.560 474.000 460.820 474.260 ;
        RECT 316.120 32.000 316.380 32.260 ;
        RECT 458.720 32.000 458.980 32.260 ;
      LAYER met2 ;
        RECT 460.810 500.000 461.090 504.000 ;
        RECT 460.850 498.340 460.990 500.000 ;
        RECT 460.620 498.200 460.990 498.340 ;
        RECT 460.620 474.290 460.760 498.200 ;
        RECT 458.720 473.970 458.980 474.290 ;
        RECT 460.560 473.970 460.820 474.290 ;
        RECT 458.780 32.290 458.920 473.970 ;
        RECT 316.120 31.970 316.380 32.290 ;
        RECT 458.720 31.970 458.980 32.290 ;
        RECT 316.180 2.400 316.320 31.970 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.140 499.500 462.460 499.760 ;
        RECT 462.230 499.080 462.370 499.500 ;
        RECT 461.910 498.880 462.370 499.080 ;
        RECT 461.910 498.820 462.230 498.880 ;
      LAYER via ;
        RECT 462.170 499.500 462.430 499.760 ;
        RECT 461.940 498.820 462.200 499.080 ;
      LAYER met2 ;
        RECT 462.190 500.000 462.470 504.000 ;
        RECT 462.230 499.790 462.370 500.000 ;
        RECT 462.170 499.470 462.430 499.790 ;
        RECT 461.940 498.965 462.200 499.110 ;
        RECT 461.930 498.595 462.210 498.965 ;
        RECT 331.290 437.395 331.570 437.765 ;
        RECT 331.360 82.870 331.500 437.395 ;
        RECT 331.360 82.730 333.800 82.870 ;
        RECT 333.660 2.400 333.800 82.730 ;
        RECT 333.450 -4.800 334.010 2.400 ;
      LAYER via2 ;
        RECT 461.930 498.640 462.210 498.920 ;
        RECT 331.290 437.440 331.570 437.720 ;
      LAYER met3 ;
        RECT 461.905 498.930 462.235 498.945 ;
        RECT 463.030 498.930 463.410 498.940 ;
        RECT 461.905 498.630 463.410 498.930 ;
        RECT 461.905 498.615 462.235 498.630 ;
        RECT 463.030 498.620 463.410 498.630 ;
        RECT 331.265 437.730 331.595 437.745 ;
        RECT 463.030 437.730 463.410 437.740 ;
        RECT 331.265 437.430 463.410 437.730 ;
        RECT 331.265 437.415 331.595 437.430 ;
        RECT 463.030 437.420 463.410 437.430 ;
      LAYER via3 ;
        RECT 463.060 498.620 463.380 498.940 ;
        RECT 463.060 437.420 463.380 437.740 ;
      LAYER met4 ;
        RECT 463.055 498.615 463.385 498.945 ;
        RECT 463.070 437.745 463.370 498.615 ;
        RECT 463.055 437.415 463.385 437.745 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 463.520 499.360 463.840 499.420 ;
        RECT 463.380 499.160 463.840 499.360 ;
        RECT 463.380 498.740 463.520 499.160 ;
        RECT 463.290 498.480 463.610 498.740 ;
      LAYER via ;
        RECT 463.550 499.160 463.810 499.420 ;
        RECT 463.320 498.480 463.580 498.740 ;
      LAYER met2 ;
        RECT 463.570 500.000 463.850 504.000 ;
        RECT 463.610 499.450 463.750 500.000 ;
        RECT 463.550 499.130 463.810 499.450 ;
        RECT 463.320 498.450 463.580 498.770 ;
        RECT 463.380 484.685 463.520 498.450 ;
        RECT 463.310 484.315 463.590 484.685 ;
        RECT 345.090 438.075 345.370 438.445 ;
        RECT 345.160 82.870 345.300 438.075 ;
        RECT 345.160 82.730 349.440 82.870 ;
        RECT 349.300 1.770 349.440 82.730 ;
        RECT 351.390 1.770 351.950 2.400 ;
        RECT 349.300 1.630 351.950 1.770 ;
        RECT 351.390 -4.800 351.950 1.630 ;
      LAYER via2 ;
        RECT 463.310 484.360 463.590 484.640 ;
        RECT 345.090 438.120 345.370 438.400 ;
      LAYER met3 ;
        RECT 463.285 484.650 463.615 484.665 ;
        RECT 463.950 484.650 464.330 484.660 ;
        RECT 463.285 484.350 464.330 484.650 ;
        RECT 463.285 484.335 463.615 484.350 ;
        RECT 463.950 484.340 464.330 484.350 ;
        RECT 345.065 438.410 345.395 438.425 ;
        RECT 463.950 438.410 464.330 438.420 ;
        RECT 345.065 438.110 464.330 438.410 ;
        RECT 345.065 438.095 345.395 438.110 ;
        RECT 463.950 438.100 464.330 438.110 ;
      LAYER via3 ;
        RECT 463.980 484.340 464.300 484.660 ;
        RECT 463.980 438.100 464.300 438.420 ;
      LAYER met4 ;
        RECT 463.975 484.335 464.305 484.665 ;
        RECT 463.990 438.425 464.290 484.335 ;
        RECT 463.975 438.095 464.305 438.425 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 466.050 472.160 466.370 472.220 ;
        RECT 468.350 472.160 468.670 472.220 ;
        RECT 466.050 472.020 468.670 472.160 ;
        RECT 466.050 471.960 466.370 472.020 ;
        RECT 468.350 471.960 468.670 472.020 ;
        RECT 368.990 33.560 369.310 33.620 ;
        RECT 468.350 33.560 468.670 33.620 ;
        RECT 368.990 33.420 468.670 33.560 ;
        RECT 368.990 33.360 369.310 33.420 ;
        RECT 468.350 33.360 468.670 33.420 ;
      LAYER via ;
        RECT 466.080 471.960 466.340 472.220 ;
        RECT 468.380 471.960 468.640 472.220 ;
        RECT 369.020 33.360 369.280 33.620 ;
        RECT 468.380 33.360 468.640 33.620 ;
      LAYER met2 ;
        RECT 464.950 500.000 465.230 504.000 ;
        RECT 464.990 499.700 465.130 500.000 ;
        RECT 464.990 499.560 465.360 499.700 ;
        RECT 465.220 487.970 465.360 499.560 ;
        RECT 465.220 487.830 465.820 487.970 ;
        RECT 465.680 473.690 465.820 487.830 ;
        RECT 465.680 473.550 466.280 473.690 ;
        RECT 466.140 472.250 466.280 473.550 ;
        RECT 466.080 471.930 466.340 472.250 ;
        RECT 468.380 471.930 468.640 472.250 ;
        RECT 468.440 33.650 468.580 471.930 ;
        RECT 369.020 33.330 369.280 33.650 ;
        RECT 468.380 33.330 468.640 33.650 ;
        RECT 369.080 2.400 369.220 33.330 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 465.130 487.460 465.450 487.520 ;
        RECT 466.510 487.460 466.830 487.520 ;
        RECT 465.130 487.320 466.830 487.460 ;
        RECT 465.130 487.260 465.450 487.320 ;
        RECT 466.510 487.260 466.830 487.320 ;
        RECT 386.930 40.360 387.250 40.420 ;
        RECT 465.130 40.360 465.450 40.420 ;
        RECT 386.930 40.220 465.450 40.360 ;
        RECT 386.930 40.160 387.250 40.220 ;
        RECT 465.130 40.160 465.450 40.220 ;
      LAYER via ;
        RECT 465.160 487.260 465.420 487.520 ;
        RECT 466.540 487.260 466.800 487.520 ;
        RECT 386.960 40.160 387.220 40.420 ;
        RECT 465.160 40.160 465.420 40.420 ;
      LAYER met2 ;
        RECT 466.330 500.000 466.610 504.000 ;
        RECT 466.370 498.680 466.510 500.000 ;
        RECT 466.370 498.540 466.740 498.680 ;
        RECT 466.600 487.550 466.740 498.540 ;
        RECT 465.160 487.230 465.420 487.550 ;
        RECT 466.540 487.230 466.800 487.550 ;
        RECT 465.220 40.450 465.360 487.230 ;
        RECT 386.960 40.130 387.220 40.450 ;
        RECT 465.160 40.130 465.420 40.450 ;
        RECT 387.020 2.400 387.160 40.130 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 467.660 499.500 467.980 499.760 ;
        RECT 467.750 498.060 467.890 499.500 ;
        RECT 467.430 497.860 467.890 498.060 ;
        RECT 467.430 497.800 467.750 497.860 ;
        RECT 464.670 472.500 464.990 472.560 ;
        RECT 467.430 472.500 467.750 472.560 ;
        RECT 464.670 472.360 467.750 472.500 ;
        RECT 464.670 472.300 464.990 472.360 ;
        RECT 467.430 472.300 467.750 472.360 ;
        RECT 404.410 40.700 404.730 40.760 ;
        RECT 464.670 40.700 464.990 40.760 ;
        RECT 404.410 40.560 464.990 40.700 ;
        RECT 404.410 40.500 404.730 40.560 ;
        RECT 464.670 40.500 464.990 40.560 ;
      LAYER via ;
        RECT 467.690 499.500 467.950 499.760 ;
        RECT 467.460 497.800 467.720 498.060 ;
        RECT 464.700 472.300 464.960 472.560 ;
        RECT 467.460 472.300 467.720 472.560 ;
        RECT 404.440 40.500 404.700 40.760 ;
        RECT 464.700 40.500 464.960 40.760 ;
      LAYER met2 ;
        RECT 467.710 500.000 467.990 504.000 ;
        RECT 467.750 499.790 467.890 500.000 ;
        RECT 467.690 499.470 467.950 499.790 ;
        RECT 467.460 497.770 467.720 498.090 ;
        RECT 467.520 472.590 467.660 497.770 ;
        RECT 464.700 472.270 464.960 472.590 ;
        RECT 467.460 472.270 467.720 472.590 ;
        RECT 464.760 40.790 464.900 472.270 ;
        RECT 404.440 40.470 404.700 40.790 ;
        RECT 464.700 40.470 464.960 40.790 ;
        RECT 404.500 2.400 404.640 40.470 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.490 500.000 441.770 504.000 ;
        RECT 441.530 498.680 441.670 500.000 ;
        RECT 441.530 498.540 441.900 498.680 ;
        RECT 441.760 488.085 441.900 498.540 ;
        RECT 441.690 487.715 441.970 488.085 ;
        RECT 67.710 23.955 67.990 24.325 ;
        RECT 67.780 2.400 67.920 23.955 ;
        RECT 67.570 -4.800 68.130 2.400 ;
      LAYER via2 ;
        RECT 441.690 487.760 441.970 488.040 ;
        RECT 67.710 24.000 67.990 24.280 ;
      LAYER met3 ;
        RECT 441.665 488.060 441.995 488.065 ;
        RECT 441.665 488.050 442.250 488.060 ;
        RECT 441.665 487.750 442.450 488.050 ;
        RECT 441.665 487.740 442.250 487.750 ;
        RECT 441.665 487.735 441.995 487.740 ;
        RECT 67.685 24.290 68.015 24.305 ;
        RECT 441.870 24.290 442.250 24.300 ;
        RECT 67.685 23.990 442.250 24.290 ;
        RECT 67.685 23.975 68.015 23.990 ;
        RECT 441.870 23.980 442.250 23.990 ;
      LAYER via3 ;
        RECT 441.900 487.740 442.220 488.060 ;
        RECT 441.900 23.980 442.220 24.300 ;
      LAYER met4 ;
        RECT 441.895 487.735 442.225 488.065 ;
        RECT 441.910 24.305 442.210 487.735 ;
        RECT 441.895 23.975 442.225 24.305 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.040 499.700 469.360 499.760 ;
        RECT 468.900 499.500 469.360 499.700 ;
        RECT 468.900 498.400 469.040 499.500 ;
        RECT 468.810 498.140 469.130 498.400 ;
      LAYER via ;
        RECT 469.070 499.500 469.330 499.760 ;
        RECT 468.840 498.140 469.100 498.400 ;
      LAYER met2 ;
        RECT 469.090 500.000 469.370 504.000 ;
        RECT 469.130 499.790 469.270 500.000 ;
        RECT 469.070 499.470 469.330 499.790 ;
        RECT 468.840 498.110 469.100 498.430 ;
        RECT 468.900 488.085 469.040 498.110 ;
        RECT 468.830 487.715 469.110 488.085 ;
        RECT 422.370 16.475 422.650 16.845 ;
        RECT 422.440 2.400 422.580 16.475 ;
        RECT 422.230 -4.800 422.790 2.400 ;
      LAYER via2 ;
        RECT 468.830 487.760 469.110 488.040 ;
        RECT 422.370 16.520 422.650 16.800 ;
      LAYER met3 ;
        RECT 468.805 488.050 469.135 488.065 ;
        RECT 470.390 488.050 470.770 488.060 ;
        RECT 468.805 487.750 470.770 488.050 ;
        RECT 468.805 487.735 469.135 487.750 ;
        RECT 470.390 487.740 470.770 487.750 ;
        RECT 422.345 16.810 422.675 16.825 ;
        RECT 470.390 16.810 470.770 16.820 ;
        RECT 422.345 16.510 470.770 16.810 ;
        RECT 422.345 16.495 422.675 16.510 ;
        RECT 470.390 16.500 470.770 16.510 ;
      LAYER via3 ;
        RECT 470.420 487.740 470.740 488.060 ;
        RECT 470.420 16.500 470.740 16.820 ;
      LAYER met4 ;
        RECT 470.415 487.735 470.745 488.065 ;
        RECT 470.430 16.825 470.730 487.735 ;
        RECT 470.415 16.495 470.745 16.825 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 470.420 499.500 470.740 499.760 ;
        RECT 470.510 498.740 470.650 499.500 ;
        RECT 470.190 498.540 470.650 498.740 ;
        RECT 470.190 498.480 470.510 498.540 ;
        RECT 437.070 482.020 437.390 482.080 ;
        RECT 470.190 482.020 470.510 482.080 ;
        RECT 437.070 481.880 470.510 482.020 ;
        RECT 437.070 481.820 437.390 481.880 ;
        RECT 470.190 481.820 470.510 481.880 ;
      LAYER via ;
        RECT 470.450 499.500 470.710 499.760 ;
        RECT 470.220 498.480 470.480 498.740 ;
        RECT 437.100 481.820 437.360 482.080 ;
        RECT 470.220 481.820 470.480 482.080 ;
      LAYER met2 ;
        RECT 470.470 500.000 470.750 504.000 ;
        RECT 470.510 499.790 470.650 500.000 ;
        RECT 470.450 499.470 470.710 499.790 ;
        RECT 470.220 498.450 470.480 498.770 ;
        RECT 470.280 482.110 470.420 498.450 ;
        RECT 437.100 481.790 437.360 482.110 ;
        RECT 470.220 481.790 470.480 482.110 ;
        RECT 437.160 2.450 437.300 481.790 ;
        RECT 437.160 2.310 437.760 2.450 ;
        RECT 437.620 1.770 437.760 2.310 ;
        RECT 439.710 1.770 440.270 2.400 ;
        RECT 437.620 1.630 440.270 1.770 ;
        RECT 439.710 -4.800 440.270 1.630 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 471.800 498.820 472.120 499.080 ;
        RECT 471.890 498.400 472.030 498.820 ;
        RECT 471.890 498.200 472.350 498.400 ;
        RECT 472.030 498.140 472.350 498.200 ;
        RECT 472.030 471.820 472.350 471.880 ;
        RECT 473.410 471.820 473.730 471.880 ;
        RECT 472.030 471.680 473.730 471.820 ;
        RECT 472.030 471.620 472.350 471.680 ;
        RECT 473.410 471.620 473.730 471.680 ;
        RECT 466.510 220.900 466.830 220.960 ;
        RECT 473.410 220.900 473.730 220.960 ;
        RECT 466.510 220.760 473.730 220.900 ;
        RECT 466.510 220.700 466.830 220.760 ;
        RECT 473.410 220.700 473.730 220.760 ;
        RECT 457.770 17.580 458.090 17.640 ;
        RECT 466.510 17.580 466.830 17.640 ;
        RECT 457.770 17.440 466.830 17.580 ;
        RECT 457.770 17.380 458.090 17.440 ;
        RECT 466.510 17.380 466.830 17.440 ;
      LAYER via ;
        RECT 471.830 498.820 472.090 499.080 ;
        RECT 472.060 498.140 472.320 498.400 ;
        RECT 472.060 471.620 472.320 471.880 ;
        RECT 473.440 471.620 473.700 471.880 ;
        RECT 466.540 220.700 466.800 220.960 ;
        RECT 473.440 220.700 473.700 220.960 ;
        RECT 457.800 17.380 458.060 17.640 ;
        RECT 466.540 17.380 466.800 17.640 ;
      LAYER met2 ;
        RECT 471.850 500.000 472.130 504.000 ;
        RECT 471.890 499.110 472.030 500.000 ;
        RECT 471.830 498.790 472.090 499.110 ;
        RECT 472.060 498.110 472.320 498.430 ;
        RECT 472.120 471.910 472.260 498.110 ;
        RECT 472.060 471.590 472.320 471.910 ;
        RECT 473.440 471.590 473.700 471.910 ;
        RECT 473.500 220.990 473.640 471.590 ;
        RECT 466.540 220.670 466.800 220.990 ;
        RECT 473.440 220.670 473.700 220.990 ;
        RECT 466.600 17.670 466.740 220.670 ;
        RECT 457.800 17.350 458.060 17.670 ;
        RECT 466.540 17.350 466.800 17.670 ;
        RECT 457.860 2.400 458.000 17.350 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.230 500.000 473.510 504.000 ;
        RECT 473.270 499.815 473.410 500.000 ;
        RECT 473.200 499.445 473.480 499.815 ;
        RECT 473.890 496.555 474.170 496.925 ;
        RECT 473.960 1.770 474.100 496.555 ;
        RECT 475.590 1.770 476.150 2.400 ;
        RECT 473.960 1.630 476.150 1.770 ;
        RECT 475.590 -4.800 476.150 1.630 ;
      LAYER via2 ;
        RECT 473.200 499.490 473.480 499.770 ;
        RECT 473.890 496.600 474.170 496.880 ;
      LAYER met3 ;
        RECT 473.175 499.465 473.505 499.795 ;
        RECT 473.190 496.890 473.490 499.465 ;
        RECT 473.865 496.890 474.195 496.905 ;
        RECT 473.190 496.590 474.195 496.890 ;
        RECT 473.865 496.575 474.195 496.590 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 474.560 498.820 474.880 499.080 ;
        RECT 474.650 497.660 474.790 498.820 ;
        RECT 474.650 497.520 475.480 497.660 ;
        RECT 471.570 496.980 471.890 497.040 ;
        RECT 475.340 496.980 475.480 497.520 ;
        RECT 471.570 496.840 475.480 496.980 ;
        RECT 471.570 496.780 471.890 496.840 ;
        RECT 471.110 15.880 471.430 15.940 ;
        RECT 493.190 15.880 493.510 15.940 ;
        RECT 471.110 15.740 493.510 15.880 ;
        RECT 471.110 15.680 471.430 15.740 ;
        RECT 493.190 15.680 493.510 15.740 ;
      LAYER via ;
        RECT 474.590 498.820 474.850 499.080 ;
        RECT 471.600 496.780 471.860 497.040 ;
        RECT 471.140 15.680 471.400 15.940 ;
        RECT 493.220 15.680 493.480 15.940 ;
      LAYER met2 ;
        RECT 474.610 500.000 474.890 504.000 ;
        RECT 474.650 499.110 474.790 500.000 ;
        RECT 474.590 498.790 474.850 499.110 ;
        RECT 471.600 496.750 471.860 497.070 ;
        RECT 471.660 468.250 471.800 496.750 ;
        RECT 471.200 468.110 471.800 468.250 ;
        RECT 471.200 15.970 471.340 468.110 ;
        RECT 471.140 15.650 471.400 15.970 ;
        RECT 493.220 15.650 493.480 15.970 ;
        RECT 493.280 2.400 493.420 15.650 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.170 471.820 476.490 471.880 ;
        RECT 478.930 471.820 479.250 471.880 ;
        RECT 476.170 471.680 479.250 471.820 ;
        RECT 476.170 471.620 476.490 471.680 ;
        RECT 478.930 471.620 479.250 471.680 ;
        RECT 478.930 20.980 479.250 21.040 ;
        RECT 511.130 20.980 511.450 21.040 ;
        RECT 478.930 20.840 511.450 20.980 ;
        RECT 478.930 20.780 479.250 20.840 ;
        RECT 511.130 20.780 511.450 20.840 ;
      LAYER via ;
        RECT 476.200 471.620 476.460 471.880 ;
        RECT 478.960 471.620 479.220 471.880 ;
        RECT 478.960 20.780 479.220 21.040 ;
        RECT 511.160 20.780 511.420 21.040 ;
      LAYER met2 ;
        RECT 475.990 500.000 476.270 504.000 ;
        RECT 476.030 499.815 476.170 500.000 ;
        RECT 475.960 499.445 476.240 499.815 ;
        RECT 475.960 498.680 476.240 498.965 ;
        RECT 475.960 498.595 476.400 498.680 ;
        RECT 476.030 498.540 476.400 498.595 ;
        RECT 476.260 471.910 476.400 498.540 ;
        RECT 476.200 471.590 476.460 471.910 ;
        RECT 478.960 471.590 479.220 471.910 ;
        RECT 479.020 21.070 479.160 471.590 ;
        RECT 478.960 20.750 479.220 21.070 ;
        RECT 511.160 20.750 511.420 21.070 ;
        RECT 511.220 2.400 511.360 20.750 ;
        RECT 511.010 -4.800 511.570 2.400 ;
      LAYER via2 ;
        RECT 475.960 499.490 476.240 499.770 ;
        RECT 475.960 498.640 476.240 498.920 ;
      LAYER met3 ;
        RECT 475.935 499.465 476.265 499.795 ;
        RECT 475.950 498.945 476.250 499.465 ;
        RECT 475.935 498.615 476.265 498.945 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 477.320 499.160 477.640 499.420 ;
        RECT 477.410 498.000 477.550 499.160 ;
        RECT 477.180 497.860 477.550 498.000 ;
        RECT 477.180 496.980 477.320 497.860 ;
        RECT 478.470 496.980 478.790 497.040 ;
        RECT 477.180 496.840 478.790 496.980 ;
        RECT 478.470 496.780 478.790 496.840 ;
        RECT 478.470 27.440 478.790 27.500 ;
        RECT 528.610 27.440 528.930 27.500 ;
        RECT 478.470 27.300 528.930 27.440 ;
        RECT 478.470 27.240 478.790 27.300 ;
        RECT 528.610 27.240 528.930 27.300 ;
      LAYER via ;
        RECT 477.350 499.160 477.610 499.420 ;
        RECT 478.500 496.780 478.760 497.040 ;
        RECT 478.500 27.240 478.760 27.500 ;
        RECT 528.640 27.240 528.900 27.500 ;
      LAYER met2 ;
        RECT 477.370 500.000 477.650 504.000 ;
        RECT 477.410 499.450 477.550 500.000 ;
        RECT 477.350 499.130 477.610 499.450 ;
        RECT 478.500 496.750 478.760 497.070 ;
        RECT 478.560 27.530 478.700 496.750 ;
        RECT 478.500 27.210 478.760 27.530 ;
        RECT 528.640 27.210 528.900 27.530 ;
        RECT 528.700 2.400 528.840 27.210 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 478.700 499.360 479.020 499.420 ;
        RECT 478.700 499.160 479.160 499.360 ;
        RECT 479.020 498.740 479.160 499.160 ;
        RECT 478.930 498.480 479.250 498.740 ;
        RECT 479.850 26.760 480.170 26.820 ;
        RECT 546.550 26.760 546.870 26.820 ;
        RECT 479.850 26.620 546.870 26.760 ;
        RECT 479.850 26.560 480.170 26.620 ;
        RECT 546.550 26.560 546.870 26.620 ;
      LAYER via ;
        RECT 478.730 499.160 478.990 499.420 ;
        RECT 478.960 498.480 479.220 498.740 ;
        RECT 479.880 26.560 480.140 26.820 ;
        RECT 546.580 26.560 546.840 26.820 ;
      LAYER met2 ;
        RECT 478.750 500.000 479.030 504.000 ;
        RECT 478.790 499.450 478.930 500.000 ;
        RECT 478.730 499.130 478.990 499.450 ;
        RECT 478.960 498.450 479.220 498.770 ;
        RECT 479.020 473.010 479.160 498.450 ;
        RECT 479.020 472.870 480.080 473.010 ;
        RECT 479.940 26.850 480.080 472.870 ;
        RECT 479.880 26.530 480.140 26.850 ;
        RECT 546.580 26.530 546.840 26.850 ;
        RECT 546.640 2.400 546.780 26.530 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 480.080 499.500 480.400 499.760 ;
        RECT 480.170 498.000 480.310 499.500 ;
        RECT 480.770 498.000 481.090 498.060 ;
        RECT 480.170 497.860 481.090 498.000 ;
        RECT 480.770 497.800 481.090 497.860 ;
        RECT 478.010 449.040 478.330 449.100 ;
        RECT 480.770 449.040 481.090 449.100 ;
        RECT 478.010 448.900 481.090 449.040 ;
        RECT 478.010 448.840 478.330 448.900 ;
        RECT 480.770 448.840 481.090 448.900 ;
        RECT 478.010 26.080 478.330 26.140 ;
        RECT 564.030 26.080 564.350 26.140 ;
        RECT 478.010 25.940 564.350 26.080 ;
        RECT 478.010 25.880 478.330 25.940 ;
        RECT 564.030 25.880 564.350 25.940 ;
      LAYER via ;
        RECT 480.110 499.500 480.370 499.760 ;
        RECT 480.800 497.800 481.060 498.060 ;
        RECT 478.040 448.840 478.300 449.100 ;
        RECT 480.800 448.840 481.060 449.100 ;
        RECT 478.040 25.880 478.300 26.140 ;
        RECT 564.060 25.880 564.320 26.140 ;
      LAYER met2 ;
        RECT 480.130 500.000 480.410 504.000 ;
        RECT 480.170 499.790 480.310 500.000 ;
        RECT 480.110 499.470 480.370 499.790 ;
        RECT 480.800 497.770 481.060 498.090 ;
        RECT 480.860 449.130 481.000 497.770 ;
        RECT 478.040 448.810 478.300 449.130 ;
        RECT 480.800 448.810 481.060 449.130 ;
        RECT 478.100 26.170 478.240 448.810 ;
        RECT 478.040 25.850 478.300 26.170 ;
        RECT 564.060 25.850 564.320 26.170 ;
        RECT 564.120 2.400 564.260 25.850 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.510 500.000 481.790 504.000 ;
        RECT 481.550 499.645 481.690 500.000 ;
        RECT 481.480 499.275 481.760 499.645 ;
        RECT 581.990 16.475 582.270 16.845 ;
        RECT 582.060 2.400 582.200 16.475 ;
        RECT 581.850 -4.800 582.410 2.400 ;
      LAYER via2 ;
        RECT 481.480 499.320 481.760 499.600 ;
        RECT 581.990 16.520 582.270 16.800 ;
      LAYER met3 ;
        RECT 480.510 499.610 480.890 499.620 ;
        RECT 481.455 499.610 481.785 499.625 ;
        RECT 480.510 499.310 481.785 499.610 ;
        RECT 480.510 499.300 480.890 499.310 ;
        RECT 481.455 499.295 481.785 499.310 ;
        RECT 480.510 16.810 480.890 16.820 ;
        RECT 581.965 16.810 582.295 16.825 ;
        RECT 480.510 16.510 582.295 16.810 ;
        RECT 480.510 16.500 480.890 16.510 ;
        RECT 581.965 16.495 582.295 16.510 ;
      LAYER via3 ;
        RECT 480.540 499.300 480.860 499.620 ;
        RECT 480.540 16.500 480.860 16.820 ;
      LAYER met4 ;
        RECT 480.535 499.295 480.865 499.625 ;
        RECT 480.550 16.825 480.850 499.295 ;
        RECT 480.535 16.495 480.865 16.825 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 91.150 38.320 91.470 38.380 ;
        RECT 444.890 38.320 445.210 38.380 ;
        RECT 91.150 38.180 445.210 38.320 ;
        RECT 91.150 38.120 91.470 38.180 ;
        RECT 444.890 38.120 445.210 38.180 ;
      LAYER via ;
        RECT 91.180 38.120 91.440 38.380 ;
        RECT 444.920 38.120 445.180 38.380 ;
      LAYER met2 ;
        RECT 443.330 500.000 443.610 504.000 ;
        RECT 443.370 499.020 443.510 500.000 ;
        RECT 443.140 498.880 443.510 499.020 ;
        RECT 443.140 498.285 443.280 498.880 ;
        RECT 443.070 497.915 443.350 498.285 ;
        RECT 444.450 497.915 444.730 498.285 ;
        RECT 444.520 491.200 444.660 497.915 ;
        RECT 444.520 491.060 445.120 491.200 ;
        RECT 444.980 38.410 445.120 491.060 ;
        RECT 91.180 38.090 91.440 38.410 ;
        RECT 444.920 38.090 445.180 38.410 ;
        RECT 91.240 2.400 91.380 38.090 ;
        RECT 91.030 -4.800 91.590 2.400 ;
      LAYER via2 ;
        RECT 443.070 497.960 443.350 498.240 ;
        RECT 444.450 497.960 444.730 498.240 ;
      LAYER met3 ;
        RECT 443.045 498.250 443.375 498.265 ;
        RECT 444.425 498.250 444.755 498.265 ;
        RECT 443.045 497.950 444.755 498.250 ;
        RECT 443.045 497.935 443.375 497.950 ;
        RECT 444.425 497.935 444.755 497.950 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 482.930 500.240 483.530 500.380 ;
        RECT 482.930 500.040 483.070 500.240 ;
        RECT 482.700 499.900 483.070 500.040 ;
        RECT 482.700 499.420 482.840 499.900 ;
        RECT 482.700 499.360 483.160 499.420 ;
        RECT 483.390 499.360 483.530 500.240 ;
        RECT 482.700 499.220 483.530 499.360 ;
        RECT 482.700 499.160 483.160 499.220 ;
        RECT 482.700 498.000 482.840 499.160 ;
        RECT 482.700 497.860 486.060 498.000 ;
        RECT 485.920 497.720 486.060 497.860 ;
        RECT 485.830 497.460 486.150 497.720 ;
        RECT 486.290 25.740 486.610 25.800 ;
        RECT 599.450 25.740 599.770 25.800 ;
        RECT 486.290 25.600 599.770 25.740 ;
        RECT 486.290 25.540 486.610 25.600 ;
        RECT 599.450 25.540 599.770 25.600 ;
      LAYER via ;
        RECT 482.870 499.160 483.130 499.420 ;
        RECT 485.860 497.460 486.120 497.720 ;
        RECT 486.320 25.540 486.580 25.800 ;
        RECT 599.480 25.540 599.740 25.800 ;
      LAYER met2 ;
        RECT 482.890 500.000 483.170 504.000 ;
        RECT 482.930 499.450 483.070 500.000 ;
        RECT 482.870 499.130 483.130 499.450 ;
        RECT 485.860 497.430 486.120 497.750 ;
        RECT 485.920 473.010 486.060 497.430 ;
        RECT 485.920 472.870 486.520 473.010 ;
        RECT 486.380 25.830 486.520 472.870 ;
        RECT 486.320 25.510 486.580 25.830 ;
        RECT 599.480 25.510 599.740 25.830 ;
        RECT 599.540 2.400 599.680 25.510 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 484.450 473.320 484.770 473.580 ;
        RECT 484.540 473.180 484.680 473.320 ;
        RECT 484.540 473.040 487.440 473.180 ;
        RECT 487.300 472.900 487.440 473.040 ;
        RECT 487.210 472.640 487.530 472.900 ;
        RECT 486.750 24.380 487.070 24.440 ;
        RECT 617.390 24.380 617.710 24.440 ;
        RECT 486.750 24.240 617.710 24.380 ;
        RECT 486.750 24.180 487.070 24.240 ;
        RECT 617.390 24.180 617.710 24.240 ;
      LAYER via ;
        RECT 484.480 473.320 484.740 473.580 ;
        RECT 487.240 472.640 487.500 472.900 ;
        RECT 486.780 24.180 487.040 24.440 ;
        RECT 617.420 24.180 617.680 24.440 ;
      LAYER met2 ;
        RECT 484.270 500.000 484.550 504.000 ;
        RECT 484.310 498.340 484.450 500.000 ;
        RECT 484.310 498.200 484.680 498.340 ;
        RECT 484.540 473.610 484.680 498.200 ;
        RECT 484.480 473.290 484.740 473.610 ;
        RECT 487.240 472.610 487.500 472.930 ;
        RECT 487.300 472.330 487.440 472.610 ;
        RECT 486.840 472.190 487.440 472.330 ;
        RECT 486.840 24.470 486.980 472.190 ;
        RECT 486.780 24.150 487.040 24.470 ;
        RECT 617.420 24.150 617.680 24.470 ;
        RECT 617.480 2.400 617.620 24.150 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 445.120 499.500 445.440 499.760 ;
        RECT 445.210 499.080 445.350 499.500 ;
        RECT 445.210 498.880 445.670 499.080 ;
        RECT 445.350 498.820 445.670 498.880 ;
        RECT 442.590 491.880 442.910 491.940 ;
        RECT 444.890 491.880 445.210 491.940 ;
        RECT 442.590 491.740 445.210 491.880 ;
        RECT 442.590 491.680 442.910 491.740 ;
        RECT 444.890 491.680 445.210 491.740 ;
        RECT 115.070 24.720 115.390 24.780 ;
        RECT 442.590 24.720 442.910 24.780 ;
        RECT 115.070 24.580 442.910 24.720 ;
        RECT 115.070 24.520 115.390 24.580 ;
        RECT 442.590 24.520 442.910 24.580 ;
      LAYER via ;
        RECT 445.150 499.500 445.410 499.760 ;
        RECT 445.380 498.820 445.640 499.080 ;
        RECT 442.620 491.680 442.880 491.940 ;
        RECT 444.920 491.680 445.180 491.940 ;
        RECT 115.100 24.520 115.360 24.780 ;
        RECT 442.620 24.520 442.880 24.780 ;
      LAYER met2 ;
        RECT 445.170 500.000 445.450 504.000 ;
        RECT 445.210 499.790 445.350 500.000 ;
        RECT 445.150 499.470 445.410 499.790 ;
        RECT 445.380 498.790 445.640 499.110 ;
        RECT 445.440 498.170 445.580 498.790 ;
        RECT 444.980 498.030 445.580 498.170 ;
        RECT 444.980 491.970 445.120 498.030 ;
        RECT 442.620 491.650 442.880 491.970 ;
        RECT 444.920 491.650 445.180 491.970 ;
        RECT 442.680 24.810 442.820 491.650 ;
        RECT 115.100 24.490 115.360 24.810 ;
        RECT 442.620 24.490 442.880 24.810 ;
        RECT 115.160 2.400 115.300 24.490 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 444.430 487.120 444.750 487.180 ;
        RECT 446.730 487.120 447.050 487.180 ;
        RECT 444.430 486.980 447.050 487.120 ;
        RECT 444.430 486.920 444.750 486.980 ;
        RECT 446.730 486.920 447.050 486.980 ;
        RECT 138.530 39.000 138.850 39.060 ;
        RECT 444.430 39.000 444.750 39.060 ;
        RECT 138.530 38.860 444.750 39.000 ;
        RECT 138.530 38.800 138.850 38.860 ;
        RECT 444.430 38.800 444.750 38.860 ;
      LAYER via ;
        RECT 444.460 486.920 444.720 487.180 ;
        RECT 446.760 486.920 447.020 487.180 ;
        RECT 138.560 38.800 138.820 39.060 ;
        RECT 444.460 38.800 444.720 39.060 ;
      LAYER met2 ;
        RECT 447.010 500.000 447.290 504.000 ;
        RECT 447.050 499.020 447.190 500.000 ;
        RECT 446.820 498.880 447.190 499.020 ;
        RECT 446.820 487.210 446.960 498.880 ;
        RECT 444.460 486.890 444.720 487.210 ;
        RECT 446.760 486.890 447.020 487.210 ;
        RECT 444.520 39.090 444.660 486.890 ;
        RECT 138.560 38.770 138.820 39.090 ;
        RECT 444.460 38.770 444.720 39.090 ;
        RECT 138.620 2.400 138.760 38.770 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.340 499.500 448.660 499.760 ;
        RECT 448.430 498.000 448.570 499.500 ;
        RECT 449.030 498.000 449.350 498.060 ;
        RECT 448.430 497.860 449.350 498.000 ;
        RECT 449.030 497.800 449.350 497.860 ;
      LAYER via ;
        RECT 448.370 499.500 448.630 499.760 ;
        RECT 449.060 497.800 449.320 498.060 ;
      LAYER met2 ;
        RECT 448.390 500.000 448.670 504.000 ;
        RECT 448.430 499.790 448.570 500.000 ;
        RECT 448.370 499.470 448.630 499.790 ;
        RECT 449.060 497.770 449.320 498.090 ;
        RECT 449.120 488.085 449.260 497.770 ;
        RECT 449.050 487.715 449.330 488.085 ;
        RECT 151.890 444.875 152.170 445.245 ;
        RECT 151.960 82.870 152.100 444.875 ;
        RECT 151.960 82.730 154.400 82.870 ;
        RECT 154.260 1.770 154.400 82.730 ;
        RECT 156.350 1.770 156.910 2.400 ;
        RECT 154.260 1.630 156.910 1.770 ;
        RECT 156.350 -4.800 156.910 1.630 ;
      LAYER via2 ;
        RECT 449.050 487.760 449.330 488.040 ;
        RECT 151.890 444.920 152.170 445.200 ;
      LAYER met3 ;
        RECT 449.025 488.060 449.355 488.065 ;
        RECT 449.025 488.050 449.610 488.060 ;
        RECT 449.025 487.750 449.810 488.050 ;
        RECT 449.025 487.740 449.610 487.750 ;
        RECT 449.025 487.735 449.355 487.740 ;
        RECT 151.865 445.210 152.195 445.225 ;
        RECT 449.230 445.210 449.610 445.220 ;
        RECT 151.865 444.910 449.610 445.210 ;
        RECT 151.865 444.895 152.195 444.910 ;
        RECT 449.230 444.900 449.610 444.910 ;
      LAYER via3 ;
        RECT 449.260 487.740 449.580 488.060 ;
        RECT 449.260 444.900 449.580 445.220 ;
      LAYER met4 ;
        RECT 449.255 487.735 449.585 488.065 ;
        RECT 449.270 445.225 449.570 487.735 ;
        RECT 449.255 444.895 449.585 445.225 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 449.720 498.820 450.040 499.080 ;
        RECT 449.810 498.060 449.950 498.820 ;
        RECT 449.490 497.860 449.950 498.060 ;
        RECT 449.490 497.800 449.810 497.860 ;
        RECT 449.490 472.500 449.810 472.560 ;
        RECT 453.170 472.500 453.490 472.560 ;
        RECT 449.490 472.360 453.490 472.500 ;
        RECT 449.490 472.300 449.810 472.360 ;
        RECT 453.170 472.300 453.490 472.360 ;
        RECT 172.570 445.300 172.890 445.360 ;
        RECT 453.170 445.300 453.490 445.360 ;
        RECT 172.570 445.160 453.490 445.300 ;
        RECT 172.570 445.100 172.890 445.160 ;
        RECT 453.170 445.100 453.490 445.160 ;
      LAYER via ;
        RECT 449.750 498.820 450.010 499.080 ;
        RECT 449.520 497.800 449.780 498.060 ;
        RECT 449.520 472.300 449.780 472.560 ;
        RECT 453.200 472.300 453.460 472.560 ;
        RECT 172.600 445.100 172.860 445.360 ;
        RECT 453.200 445.100 453.460 445.360 ;
      LAYER met2 ;
        RECT 449.770 500.000 450.050 504.000 ;
        RECT 449.810 499.110 449.950 500.000 ;
        RECT 449.750 498.790 450.010 499.110 ;
        RECT 449.520 497.770 449.780 498.090 ;
        RECT 449.580 472.590 449.720 497.770 ;
        RECT 449.520 472.270 449.780 472.590 ;
        RECT 453.200 472.270 453.460 472.590 ;
        RECT 453.260 445.390 453.400 472.270 ;
        RECT 172.600 445.070 172.860 445.390 ;
        RECT 453.200 445.070 453.460 445.390 ;
        RECT 172.660 1.770 172.800 445.070 ;
        RECT 173.830 1.770 174.390 2.400 ;
        RECT 172.660 1.630 174.390 1.770 ;
        RECT 173.830 -4.800 174.390 1.630 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 451.100 499.160 451.420 499.420 ;
        RECT 451.190 498.060 451.330 499.160 ;
        RECT 451.190 497.860 451.650 498.060 ;
        RECT 451.330 497.800 451.650 497.860 ;
        RECT 451.330 488.820 451.650 488.880 ;
        RECT 451.330 488.680 454.320 488.820 ;
        RECT 451.330 488.620 451.650 488.680 ;
        RECT 454.180 488.540 454.320 488.680 ;
        RECT 454.090 488.280 454.410 488.540 ;
        RECT 191.890 26.080 192.210 26.140 ;
        RECT 453.630 26.080 453.950 26.140 ;
        RECT 191.890 25.940 453.950 26.080 ;
        RECT 191.890 25.880 192.210 25.940 ;
        RECT 453.630 25.880 453.950 25.940 ;
      LAYER via ;
        RECT 451.130 499.160 451.390 499.420 ;
        RECT 451.360 497.800 451.620 498.060 ;
        RECT 451.360 488.620 451.620 488.880 ;
        RECT 454.120 488.280 454.380 488.540 ;
        RECT 191.920 25.880 192.180 26.140 ;
        RECT 453.660 25.880 453.920 26.140 ;
      LAYER met2 ;
        RECT 451.150 500.000 451.430 504.000 ;
        RECT 451.190 499.450 451.330 500.000 ;
        RECT 451.130 499.130 451.390 499.450 ;
        RECT 451.360 497.770 451.620 498.090 ;
        RECT 451.420 488.910 451.560 497.770 ;
        RECT 451.360 488.590 451.620 488.910 ;
        RECT 454.120 488.250 454.380 488.570 ;
        RECT 454.180 420.970 454.320 488.250 ;
        RECT 453.720 420.830 454.320 420.970 ;
        RECT 453.720 26.170 453.860 420.830 ;
        RECT 191.920 25.850 192.180 26.170 ;
        RECT 453.660 25.850 453.920 26.170 ;
        RECT 191.980 2.400 192.120 25.850 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 209.370 40.020 209.690 40.080 ;
        RECT 451.330 40.020 451.650 40.080 ;
        RECT 209.370 39.880 451.650 40.020 ;
        RECT 209.370 39.820 209.690 39.880 ;
        RECT 451.330 39.820 451.650 39.880 ;
      LAYER via ;
        RECT 209.400 39.820 209.660 40.080 ;
        RECT 451.360 39.820 451.620 40.080 ;
      LAYER met2 ;
        RECT 452.530 500.000 452.810 504.000 ;
        RECT 452.570 497.660 452.710 500.000 ;
        RECT 452.340 497.520 452.710 497.660 ;
        RECT 452.340 476.170 452.480 497.520 ;
        RECT 451.880 476.030 452.480 476.170 ;
        RECT 451.880 472.330 452.020 476.030 ;
        RECT 451.420 472.190 452.020 472.330 ;
        RECT 451.420 40.110 451.560 472.190 ;
        RECT 209.400 39.790 209.660 40.110 ;
        RECT 451.360 39.790 451.620 40.110 ;
        RECT 209.460 2.400 209.600 39.790 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 453.860 499.500 454.180 499.760 ;
        RECT 453.950 499.080 454.090 499.500 ;
        RECT 453.950 498.880 454.410 499.080 ;
        RECT 454.090 498.820 454.410 498.880 ;
        RECT 449.490 471.820 449.810 471.880 ;
        RECT 454.550 471.820 454.870 471.880 ;
        RECT 449.490 471.680 454.870 471.820 ;
        RECT 449.490 471.620 449.810 471.680 ;
        RECT 454.550 471.620 454.870 471.680 ;
        RECT 227.310 27.100 227.630 27.160 ;
        RECT 449.490 27.100 449.810 27.160 ;
        RECT 227.310 26.960 449.810 27.100 ;
        RECT 227.310 26.900 227.630 26.960 ;
        RECT 449.490 26.900 449.810 26.960 ;
      LAYER via ;
        RECT 453.890 499.500 454.150 499.760 ;
        RECT 454.120 498.820 454.380 499.080 ;
        RECT 449.520 471.620 449.780 471.880 ;
        RECT 454.580 471.620 454.840 471.880 ;
        RECT 227.340 26.900 227.600 27.160 ;
        RECT 449.520 26.900 449.780 27.160 ;
      LAYER met2 ;
        RECT 453.910 500.000 454.190 504.000 ;
        RECT 453.950 499.790 454.090 500.000 ;
        RECT 453.890 499.470 454.150 499.790 ;
        RECT 454.120 498.790 454.380 499.110 ;
        RECT 454.180 489.160 454.320 498.790 ;
        RECT 454.180 489.020 454.780 489.160 ;
        RECT 454.640 471.910 454.780 489.020 ;
        RECT 449.520 471.590 449.780 471.910 ;
        RECT 454.580 471.590 454.840 471.910 ;
        RECT 449.580 27.190 449.720 471.590 ;
        RECT 227.340 26.870 227.600 27.190 ;
        RECT 449.520 26.870 449.780 27.190 ;
        RECT 227.400 2.400 227.540 26.870 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 438.450 484.060 438.770 484.120 ;
        RECT 440.290 484.060 440.610 484.120 ;
        RECT 438.450 483.920 440.610 484.060 ;
        RECT 438.450 483.860 438.770 483.920 ;
        RECT 440.290 483.860 440.610 483.920 ;
        RECT 49.750 44.780 50.070 44.840 ;
        RECT 438.450 44.780 438.770 44.840 ;
        RECT 49.750 44.640 438.770 44.780 ;
        RECT 49.750 44.580 50.070 44.640 ;
        RECT 438.450 44.580 438.770 44.640 ;
      LAYER via ;
        RECT 438.480 483.860 438.740 484.120 ;
        RECT 440.320 483.860 440.580 484.120 ;
        RECT 49.780 44.580 50.040 44.840 ;
        RECT 438.480 44.580 438.740 44.840 ;
      LAYER met2 ;
        RECT 440.110 500.000 440.390 504.000 ;
        RECT 440.150 498.340 440.290 500.000 ;
        RECT 440.150 498.200 440.520 498.340 ;
        RECT 440.380 484.150 440.520 498.200 ;
        RECT 438.480 483.830 438.740 484.150 ;
        RECT 440.320 483.830 440.580 484.150 ;
        RECT 438.540 44.870 438.680 483.830 ;
        RECT 49.780 44.550 50.040 44.870 ;
        RECT 438.480 44.550 438.740 44.870 ;
        RECT 49.840 2.400 49.980 44.550 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.750 500.000 456.030 504.000 ;
        RECT 455.790 498.965 455.930 500.000 ;
        RECT 455.720 498.595 456.000 498.965 ;
        RECT 250.790 25.995 251.070 26.365 ;
        RECT 250.860 2.400 251.000 25.995 ;
        RECT 250.650 -4.800 251.210 2.400 ;
      LAYER via2 ;
        RECT 455.720 498.640 456.000 498.920 ;
        RECT 250.790 26.040 251.070 26.320 ;
      LAYER met3 ;
        RECT 455.695 498.940 456.025 498.945 ;
        RECT 455.670 498.930 456.050 498.940 ;
        RECT 455.240 498.630 456.050 498.930 ;
        RECT 455.670 498.620 456.050 498.630 ;
        RECT 455.695 498.615 456.025 498.620 ;
        RECT 250.765 26.330 251.095 26.345 ;
        RECT 455.670 26.330 456.050 26.340 ;
        RECT 250.765 26.030 456.050 26.330 ;
        RECT 250.765 26.015 251.095 26.030 ;
        RECT 455.670 26.020 456.050 26.030 ;
      LAYER via3 ;
        RECT 455.700 498.620 456.020 498.940 ;
        RECT 455.700 26.020 456.020 26.340 ;
      LAYER met4 ;
        RECT 455.695 498.615 456.025 498.945 ;
        RECT 455.710 26.345 456.010 498.615 ;
        RECT 455.695 26.015 456.025 26.345 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 434.770 501.060 435.090 501.120 ;
        RECT 457.080 501.060 457.400 501.120 ;
        RECT 434.770 500.920 457.400 501.060 ;
        RECT 434.770 500.860 435.090 500.920 ;
        RECT 457.080 500.860 457.400 500.920 ;
        RECT 434.770 484.740 435.090 484.800 ;
        RECT 438.910 484.740 439.230 484.800 ;
        RECT 434.770 484.600 439.230 484.740 ;
        RECT 434.770 484.540 435.090 484.600 ;
        RECT 438.910 484.540 439.230 484.600 ;
        RECT 262.270 445.640 262.590 445.700 ;
        RECT 438.910 445.640 439.230 445.700 ;
        RECT 262.270 445.500 439.230 445.640 ;
        RECT 262.270 445.440 262.590 445.500 ;
        RECT 438.910 445.440 439.230 445.500 ;
      LAYER via ;
        RECT 434.800 500.860 435.060 501.120 ;
        RECT 457.110 500.860 457.370 501.120 ;
        RECT 434.800 484.540 435.060 484.800 ;
        RECT 438.940 484.540 439.200 484.800 ;
        RECT 262.300 445.440 262.560 445.700 ;
        RECT 438.940 445.440 439.200 445.700 ;
      LAYER met2 ;
        RECT 457.130 501.150 457.410 504.000 ;
        RECT 434.800 500.830 435.060 501.150 ;
        RECT 457.110 500.830 457.410 501.150 ;
        RECT 434.860 484.830 435.000 500.830 ;
        RECT 457.130 500.000 457.410 500.830 ;
        RECT 434.800 484.510 435.060 484.830 ;
        RECT 438.940 484.510 439.200 484.830 ;
        RECT 439.000 445.730 439.140 484.510 ;
        RECT 262.300 445.410 262.560 445.730 ;
        RECT 438.940 445.410 439.200 445.730 ;
        RECT 262.360 82.870 262.500 445.410 ;
        RECT 262.360 82.730 266.640 82.870 ;
        RECT 266.500 1.770 266.640 82.730 ;
        RECT 268.590 1.770 269.150 2.400 ;
        RECT 266.500 1.630 269.150 1.770 ;
        RECT 268.590 -4.800 269.150 1.630 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 286.190 31.520 286.510 31.580 ;
        RECT 458.230 31.520 458.550 31.580 ;
        RECT 286.190 31.380 458.550 31.520 ;
        RECT 286.190 31.320 286.510 31.380 ;
        RECT 458.230 31.320 458.550 31.380 ;
      LAYER via ;
        RECT 286.220 31.320 286.480 31.580 ;
        RECT 458.260 31.320 458.520 31.580 ;
      LAYER met2 ;
        RECT 458.510 500.000 458.790 504.000 ;
        RECT 458.550 498.340 458.690 500.000 ;
        RECT 458.320 498.200 458.690 498.340 ;
        RECT 458.320 31.610 458.460 498.200 ;
        RECT 286.220 31.290 286.480 31.610 ;
        RECT 458.260 31.290 458.520 31.610 ;
        RECT 286.280 2.400 286.420 31.290 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 431.090 489.500 431.410 489.560 ;
        RECT 459.610 489.500 459.930 489.560 ;
        RECT 431.090 489.360 459.930 489.500 ;
        RECT 431.090 489.300 431.410 489.360 ;
        RECT 459.610 489.300 459.930 489.360 ;
        RECT 304.130 32.880 304.450 32.940 ;
        RECT 431.090 32.880 431.410 32.940 ;
        RECT 304.130 32.740 431.410 32.880 ;
        RECT 304.130 32.680 304.450 32.740 ;
        RECT 431.090 32.680 431.410 32.740 ;
      LAYER via ;
        RECT 431.120 489.300 431.380 489.560 ;
        RECT 459.640 489.300 459.900 489.560 ;
        RECT 304.160 32.680 304.420 32.940 ;
        RECT 431.120 32.680 431.380 32.940 ;
      LAYER met2 ;
        RECT 459.890 500.000 460.170 504.000 ;
        RECT 459.930 498.170 460.070 500.000 ;
        RECT 459.700 498.030 460.070 498.170 ;
        RECT 459.700 489.590 459.840 498.030 ;
        RECT 431.120 489.270 431.380 489.590 ;
        RECT 459.640 489.270 459.900 489.590 ;
        RECT 431.180 32.970 431.320 489.270 ;
        RECT 304.160 32.650 304.420 32.970 ;
        RECT 431.120 32.650 431.380 32.970 ;
        RECT 304.220 2.400 304.360 32.650 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.790 499.900 461.450 500.040 ;
        RECT 455.790 499.020 455.930 499.900 ;
        RECT 461.310 499.760 461.450 499.900 ;
        RECT 461.220 499.500 461.540 499.760 ;
        RECT 455.560 498.880 455.930 499.020 ;
        RECT 455.560 498.400 455.700 498.880 ;
        RECT 455.470 498.140 455.790 498.400 ;
        RECT 452.250 471.140 452.570 471.200 ;
        RECT 455.470 471.140 455.790 471.200 ;
        RECT 452.250 471.000 455.790 471.140 ;
        RECT 452.250 470.940 452.570 471.000 ;
        RECT 455.470 470.940 455.790 471.000 ;
        RECT 321.610 32.540 321.930 32.600 ;
        RECT 452.250 32.540 452.570 32.600 ;
        RECT 321.610 32.400 452.570 32.540 ;
        RECT 321.610 32.340 321.930 32.400 ;
        RECT 452.250 32.340 452.570 32.400 ;
      LAYER via ;
        RECT 461.250 499.500 461.510 499.760 ;
        RECT 455.500 498.140 455.760 498.400 ;
        RECT 452.280 470.940 452.540 471.200 ;
        RECT 455.500 470.940 455.760 471.200 ;
        RECT 321.640 32.340 321.900 32.600 ;
        RECT 452.280 32.340 452.540 32.600 ;
      LAYER met2 ;
        RECT 461.270 500.000 461.550 504.000 ;
        RECT 461.310 499.790 461.450 500.000 ;
        RECT 461.250 499.470 461.510 499.790 ;
        RECT 455.500 498.110 455.760 498.430 ;
        RECT 455.560 471.230 455.700 498.110 ;
        RECT 452.280 470.910 452.540 471.230 ;
        RECT 455.500 470.910 455.760 471.230 ;
        RECT 452.340 32.630 452.480 470.910 ;
        RECT 321.640 32.310 321.900 32.630 ;
        RECT 452.280 32.310 452.540 32.630 ;
        RECT 321.700 2.400 321.840 32.310 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.600 499.160 462.920 499.420 ;
        RECT 462.690 498.740 462.830 499.160 ;
        RECT 462.370 498.540 462.830 498.740 ;
        RECT 462.370 498.480 462.690 498.540 ;
        RECT 431.550 477.600 431.870 477.660 ;
        RECT 462.370 477.600 462.690 477.660 ;
        RECT 431.550 477.460 462.690 477.600 ;
        RECT 431.550 477.400 431.870 477.460 ;
        RECT 462.370 477.400 462.690 477.460 ;
        RECT 339.550 33.900 339.870 33.960 ;
        RECT 431.550 33.900 431.870 33.960 ;
        RECT 339.550 33.760 431.870 33.900 ;
        RECT 339.550 33.700 339.870 33.760 ;
        RECT 431.550 33.700 431.870 33.760 ;
      LAYER via ;
        RECT 462.630 499.160 462.890 499.420 ;
        RECT 462.400 498.480 462.660 498.740 ;
        RECT 431.580 477.400 431.840 477.660 ;
        RECT 462.400 477.400 462.660 477.660 ;
        RECT 339.580 33.700 339.840 33.960 ;
        RECT 431.580 33.700 431.840 33.960 ;
      LAYER met2 ;
        RECT 462.650 500.000 462.930 504.000 ;
        RECT 462.690 499.450 462.830 500.000 ;
        RECT 462.630 499.130 462.890 499.450 ;
        RECT 462.400 498.450 462.660 498.770 ;
        RECT 462.460 477.690 462.600 498.450 ;
        RECT 431.580 477.370 431.840 477.690 ;
        RECT 462.400 477.370 462.660 477.690 ;
        RECT 431.640 33.990 431.780 477.370 ;
        RECT 339.580 33.670 339.840 33.990 ;
        RECT 431.580 33.670 431.840 33.990 ;
        RECT 339.640 2.400 339.780 33.670 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 357.490 33.220 357.810 33.280 ;
        RECT 463.750 33.220 464.070 33.280 ;
        RECT 357.490 33.080 464.070 33.220 ;
        RECT 357.490 33.020 357.810 33.080 ;
        RECT 463.750 33.020 464.070 33.080 ;
      LAYER via ;
        RECT 357.520 33.020 357.780 33.280 ;
        RECT 463.780 33.020 464.040 33.280 ;
      LAYER met2 ;
        RECT 464.030 500.000 464.310 504.000 ;
        RECT 464.070 499.020 464.210 500.000 ;
        RECT 464.070 498.880 464.440 499.020 ;
        RECT 464.300 498.000 464.440 498.880 ;
        RECT 463.840 497.860 464.440 498.000 ;
        RECT 463.840 33.310 463.980 497.860 ;
        RECT 357.520 32.990 357.780 33.310 ;
        RECT 463.780 32.990 464.040 33.310 ;
        RECT 357.580 2.400 357.720 32.990 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 432.470 500.720 432.790 500.780 ;
        RECT 465.360 500.720 465.680 500.780 ;
        RECT 432.470 500.580 465.680 500.720 ;
        RECT 432.470 500.520 432.790 500.580 ;
        RECT 465.360 500.520 465.680 500.580 ;
        RECT 374.970 41.040 375.290 41.100 ;
        RECT 432.470 41.040 432.790 41.100 ;
        RECT 374.970 40.900 432.790 41.040 ;
        RECT 374.970 40.840 375.290 40.900 ;
        RECT 432.470 40.840 432.790 40.900 ;
      LAYER via ;
        RECT 432.500 500.520 432.760 500.780 ;
        RECT 465.390 500.520 465.650 500.780 ;
        RECT 375.000 40.840 375.260 41.100 ;
        RECT 432.500 40.840 432.760 41.100 ;
      LAYER met2 ;
        RECT 465.410 500.810 465.690 504.000 ;
        RECT 432.500 500.490 432.760 500.810 ;
        RECT 465.390 500.490 465.690 500.810 ;
        RECT 432.560 41.130 432.700 500.490 ;
        RECT 465.410 500.000 465.690 500.490 ;
        RECT 375.000 40.810 375.260 41.130 ;
        RECT 432.500 40.810 432.760 41.130 ;
        RECT 375.060 2.400 375.200 40.810 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 466.740 499.500 467.060 499.760 ;
        RECT 464.670 496.980 464.990 497.040 ;
        RECT 466.830 496.980 466.970 499.500 ;
        RECT 464.670 496.840 466.970 496.980 ;
        RECT 464.670 496.780 464.990 496.840 ;
        RECT 392.910 30.500 393.230 30.560 ;
        RECT 464.210 30.500 464.530 30.560 ;
        RECT 392.910 30.360 464.530 30.500 ;
        RECT 392.910 30.300 393.230 30.360 ;
        RECT 464.210 30.300 464.530 30.360 ;
      LAYER via ;
        RECT 466.770 499.500 467.030 499.760 ;
        RECT 464.700 496.780 464.960 497.040 ;
        RECT 392.940 30.300 393.200 30.560 ;
        RECT 464.240 30.300 464.500 30.560 ;
      LAYER met2 ;
        RECT 466.790 500.000 467.070 504.000 ;
        RECT 466.830 499.790 466.970 500.000 ;
        RECT 466.770 499.470 467.030 499.790 ;
        RECT 464.700 496.750 464.960 497.070 ;
        RECT 464.760 473.010 464.900 496.750 ;
        RECT 464.300 472.870 464.900 473.010 ;
        RECT 464.300 30.590 464.440 472.870 ;
        RECT 392.940 30.270 393.200 30.590 ;
        RECT 464.240 30.270 464.500 30.590 ;
        RECT 393.000 2.400 393.140 30.270 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 432.010 500.380 432.330 500.440 ;
        RECT 432.010 500.240 468.350 500.380 ;
        RECT 432.010 500.180 432.330 500.240 ;
        RECT 468.210 499.760 468.350 500.240 ;
        RECT 468.120 499.500 468.440 499.760 ;
        RECT 410.390 34.580 410.710 34.640 ;
        RECT 432.010 34.580 432.330 34.640 ;
        RECT 410.390 34.440 432.330 34.580 ;
        RECT 410.390 34.380 410.710 34.440 ;
        RECT 432.010 34.380 432.330 34.440 ;
      LAYER via ;
        RECT 432.040 500.180 432.300 500.440 ;
        RECT 468.150 499.500 468.410 499.760 ;
        RECT 410.420 34.380 410.680 34.640 ;
        RECT 432.040 34.380 432.300 34.640 ;
      LAYER met2 ;
        RECT 432.040 500.150 432.300 500.470 ;
        RECT 432.100 34.670 432.240 500.150 ;
        RECT 468.170 500.000 468.450 504.000 ;
        RECT 468.210 499.790 468.350 500.000 ;
        RECT 468.150 499.470 468.410 499.790 ;
        RECT 410.420 34.350 410.680 34.670 ;
        RECT 432.040 34.350 432.300 34.670 ;
        RECT 410.480 2.400 410.620 34.350 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 432.930 485.760 433.250 485.820 ;
        RECT 435.230 485.760 435.550 485.820 ;
        RECT 432.930 485.620 435.550 485.760 ;
        RECT 432.930 485.560 433.250 485.620 ;
        RECT 435.230 485.560 435.550 485.620 ;
        RECT 69.070 444.960 69.390 445.020 ;
        RECT 432.930 444.960 433.250 445.020 ;
        RECT 69.070 444.820 433.250 444.960 ;
        RECT 69.070 444.760 69.390 444.820 ;
        RECT 432.930 444.760 433.250 444.820 ;
      LAYER via ;
        RECT 432.960 485.560 433.220 485.820 ;
        RECT 435.260 485.560 435.520 485.820 ;
        RECT 69.100 444.760 69.360 445.020 ;
        RECT 432.960 444.760 433.220 445.020 ;
      LAYER met2 ;
        RECT 441.950 500.000 442.230 504.000 ;
        RECT 441.990 499.815 442.130 500.000 ;
        RECT 441.920 499.445 442.200 499.815 ;
        RECT 435.250 498.595 435.530 498.965 ;
        RECT 435.320 485.850 435.460 498.595 ;
        RECT 432.960 485.530 433.220 485.850 ;
        RECT 435.260 485.530 435.520 485.850 ;
        RECT 433.020 445.050 433.160 485.530 ;
        RECT 69.100 444.730 69.360 445.050 ;
        RECT 432.960 444.730 433.220 445.050 ;
        RECT 69.160 82.870 69.300 444.730 ;
        RECT 69.160 82.730 71.600 82.870 ;
        RECT 71.460 1.770 71.600 82.730 ;
        RECT 73.550 1.770 74.110 2.400 ;
        RECT 71.460 1.630 74.110 1.770 ;
        RECT 73.550 -4.800 74.110 1.630 ;
      LAYER via2 ;
        RECT 441.920 499.490 442.200 499.770 ;
        RECT 435.250 498.640 435.530 498.920 ;
      LAYER met3 ;
        RECT 441.895 499.610 442.225 499.795 ;
        RECT 440.990 499.465 442.225 499.610 ;
        RECT 440.990 499.310 442.210 499.465 ;
        RECT 435.225 498.930 435.555 498.945 ;
        RECT 440.990 498.930 441.290 499.310 ;
        RECT 435.225 498.630 441.290 498.930 ;
        RECT 435.225 498.615 435.555 498.630 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.500 499.500 469.820 499.760 ;
        RECT 469.590 499.360 469.730 499.500 ;
        RECT 469.360 499.220 469.730 499.360 ;
        RECT 469.360 497.720 469.500 499.220 ;
        RECT 469.270 497.460 469.590 497.720 ;
      LAYER via ;
        RECT 469.530 499.500 469.790 499.760 ;
        RECT 469.300 497.460 469.560 497.720 ;
      LAYER met2 ;
        RECT 469.550 500.000 469.830 504.000 ;
        RECT 469.590 499.790 469.730 500.000 ;
        RECT 469.530 499.470 469.790 499.790 ;
        RECT 469.300 497.430 469.560 497.750 ;
        RECT 469.360 488.765 469.500 497.430 ;
        RECT 469.290 488.395 469.570 488.765 ;
        RECT 428.350 17.155 428.630 17.525 ;
        RECT 428.420 2.400 428.560 17.155 ;
        RECT 428.210 -4.800 428.770 2.400 ;
      LAYER via2 ;
        RECT 469.290 488.440 469.570 488.720 ;
        RECT 428.350 17.200 428.630 17.480 ;
      LAYER met3 ;
        RECT 469.265 488.740 469.595 488.745 ;
        RECT 469.265 488.730 469.850 488.740 ;
        RECT 469.265 488.430 470.050 488.730 ;
        RECT 469.265 488.420 469.850 488.430 ;
        RECT 469.265 488.415 469.595 488.420 ;
        RECT 428.325 17.490 428.655 17.505 ;
        RECT 469.470 17.490 469.850 17.500 ;
        RECT 428.325 17.190 469.850 17.490 ;
        RECT 428.325 17.175 428.655 17.190 ;
        RECT 469.470 17.180 469.850 17.190 ;
      LAYER via3 ;
        RECT 469.500 488.420 469.820 488.740 ;
        RECT 469.500 17.180 469.820 17.500 ;
      LAYER met4 ;
        RECT 469.495 488.415 469.825 488.745 ;
        RECT 469.510 17.505 469.810 488.415 ;
        RECT 469.495 17.175 469.825 17.505 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 470.880 499.160 471.200 499.420 ;
        RECT 470.970 498.400 471.110 499.160 ;
        RECT 470.650 498.200 471.110 498.400 ;
        RECT 470.650 498.140 470.970 498.200 ;
        RECT 445.810 14.860 446.130 14.920 ;
        RECT 470.650 14.860 470.970 14.920 ;
        RECT 445.810 14.720 470.970 14.860 ;
        RECT 445.810 14.660 446.130 14.720 ;
        RECT 470.650 14.660 470.970 14.720 ;
      LAYER via ;
        RECT 470.910 499.160 471.170 499.420 ;
        RECT 470.680 498.140 470.940 498.400 ;
        RECT 445.840 14.660 446.100 14.920 ;
        RECT 470.680 14.660 470.940 14.920 ;
      LAYER met2 ;
        RECT 470.930 500.000 471.210 504.000 ;
        RECT 470.970 499.450 471.110 500.000 ;
        RECT 470.910 499.130 471.170 499.450 ;
        RECT 470.680 498.110 470.940 498.430 ;
        RECT 470.740 14.950 470.880 498.110 ;
        RECT 445.840 14.630 446.100 14.950 ;
        RECT 470.680 14.630 470.940 14.950 ;
        RECT 445.900 2.400 446.040 14.630 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 472.260 499.500 472.580 499.760 ;
        RECT 472.350 498.680 472.490 499.500 ;
        RECT 472.350 498.540 472.720 498.680 ;
        RECT 472.580 498.060 472.720 498.540 ;
        RECT 472.490 497.800 472.810 498.060 ;
        RECT 463.750 18.600 464.070 18.660 ;
        RECT 472.950 18.600 473.270 18.660 ;
        RECT 463.750 18.460 473.270 18.600 ;
        RECT 463.750 18.400 464.070 18.460 ;
        RECT 472.950 18.400 473.270 18.460 ;
      LAYER via ;
        RECT 472.290 499.500 472.550 499.760 ;
        RECT 472.520 497.800 472.780 498.060 ;
        RECT 463.780 18.400 464.040 18.660 ;
        RECT 472.980 18.400 473.240 18.660 ;
      LAYER met2 ;
        RECT 472.310 500.000 472.590 504.000 ;
        RECT 472.350 499.790 472.490 500.000 ;
        RECT 472.290 499.470 472.550 499.790 ;
        RECT 472.520 497.770 472.780 498.090 ;
        RECT 472.580 473.010 472.720 497.770 ;
        RECT 472.580 472.870 473.180 473.010 ;
        RECT 473.040 18.690 473.180 472.870 ;
        RECT 463.780 18.370 464.040 18.690 ;
        RECT 472.980 18.370 473.240 18.690 ;
        RECT 463.840 2.400 463.980 18.370 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 473.640 499.160 473.960 499.420 ;
        RECT 473.730 497.720 473.870 499.160 ;
        RECT 473.410 497.520 473.870 497.720 ;
        RECT 473.410 497.460 473.730 497.520 ;
        RECT 472.490 472.500 472.810 472.560 ;
        RECT 473.410 472.500 473.730 472.560 ;
        RECT 472.490 472.360 473.730 472.500 ;
        RECT 472.490 472.300 472.810 472.360 ;
        RECT 473.410 472.300 473.730 472.360 ;
        RECT 472.490 17.240 472.810 17.300 ;
        RECT 481.230 17.240 481.550 17.300 ;
        RECT 472.490 17.100 481.550 17.240 ;
        RECT 472.490 17.040 472.810 17.100 ;
        RECT 481.230 17.040 481.550 17.100 ;
      LAYER via ;
        RECT 473.670 499.160 473.930 499.420 ;
        RECT 473.440 497.460 473.700 497.720 ;
        RECT 472.520 472.300 472.780 472.560 ;
        RECT 473.440 472.300 473.700 472.560 ;
        RECT 472.520 17.040 472.780 17.300 ;
        RECT 481.260 17.040 481.520 17.300 ;
      LAYER met2 ;
        RECT 473.690 500.000 473.970 504.000 ;
        RECT 473.730 499.450 473.870 500.000 ;
        RECT 473.670 499.130 473.930 499.450 ;
        RECT 473.440 497.430 473.700 497.750 ;
        RECT 473.500 476.170 473.640 497.430 ;
        RECT 473.040 476.030 473.640 476.170 ;
        RECT 473.040 473.690 473.180 476.030 ;
        RECT 473.040 473.550 473.640 473.690 ;
        RECT 473.500 472.590 473.640 473.550 ;
        RECT 472.520 472.270 472.780 472.590 ;
        RECT 473.440 472.270 473.700 472.590 ;
        RECT 472.580 17.330 472.720 472.270 ;
        RECT 472.520 17.010 472.780 17.330 ;
        RECT 481.260 17.010 481.520 17.330 ;
        RECT 481.320 2.400 481.460 17.010 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 475.020 499.500 475.340 499.760 ;
        RECT 475.110 498.060 475.250 499.500 ;
        RECT 475.110 497.860 475.570 498.060 ;
        RECT 475.250 497.800 475.570 497.860 ;
        RECT 472.030 460.600 472.350 460.660 ;
        RECT 475.250 460.600 475.570 460.660 ;
        RECT 472.030 460.460 475.570 460.600 ;
        RECT 472.030 460.400 472.350 460.460 ;
        RECT 475.250 460.400 475.570 460.460 ;
        RECT 472.030 58.720 472.350 58.780 ;
        RECT 473.410 58.720 473.730 58.780 ;
        RECT 472.030 58.580 473.730 58.720 ;
        RECT 472.030 58.520 472.350 58.580 ;
        RECT 473.410 58.520 473.730 58.580 ;
        RECT 473.410 17.920 473.730 17.980 ;
        RECT 499.170 17.920 499.490 17.980 ;
        RECT 473.410 17.780 499.490 17.920 ;
        RECT 473.410 17.720 473.730 17.780 ;
        RECT 499.170 17.720 499.490 17.780 ;
      LAYER via ;
        RECT 475.050 499.500 475.310 499.760 ;
        RECT 475.280 497.800 475.540 498.060 ;
        RECT 472.060 460.400 472.320 460.660 ;
        RECT 475.280 460.400 475.540 460.660 ;
        RECT 472.060 58.520 472.320 58.780 ;
        RECT 473.440 58.520 473.700 58.780 ;
        RECT 473.440 17.720 473.700 17.980 ;
        RECT 499.200 17.720 499.460 17.980 ;
      LAYER met2 ;
        RECT 475.070 500.000 475.350 504.000 ;
        RECT 475.110 499.790 475.250 500.000 ;
        RECT 475.050 499.470 475.310 499.790 ;
        RECT 475.280 497.770 475.540 498.090 ;
        RECT 475.340 460.690 475.480 497.770 ;
        RECT 472.060 460.370 472.320 460.690 ;
        RECT 475.280 460.370 475.540 460.690 ;
        RECT 472.120 58.810 472.260 460.370 ;
        RECT 472.060 58.490 472.320 58.810 ;
        RECT 473.440 58.490 473.700 58.810 ;
        RECT 473.500 18.010 473.640 58.490 ;
        RECT 473.440 17.690 473.700 18.010 ;
        RECT 499.200 17.690 499.460 18.010 ;
        RECT 499.260 2.400 499.400 17.690 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.400 499.360 476.720 499.420 ;
        RECT 476.400 499.160 476.860 499.360 ;
        RECT 476.720 498.740 476.860 499.160 ;
        RECT 476.630 498.480 476.950 498.740 ;
        RECT 476.630 15.540 476.950 15.600 ;
        RECT 516.650 15.540 516.970 15.600 ;
        RECT 476.630 15.400 516.970 15.540 ;
        RECT 476.630 15.340 476.950 15.400 ;
        RECT 516.650 15.340 516.970 15.400 ;
      LAYER via ;
        RECT 476.430 499.160 476.690 499.420 ;
        RECT 476.660 498.480 476.920 498.740 ;
        RECT 476.660 15.340 476.920 15.600 ;
        RECT 516.680 15.340 516.940 15.600 ;
      LAYER met2 ;
        RECT 476.450 500.000 476.730 504.000 ;
        RECT 476.490 499.450 476.630 500.000 ;
        RECT 476.430 499.130 476.690 499.450 ;
        RECT 476.660 498.450 476.920 498.770 ;
        RECT 476.720 15.630 476.860 498.450 ;
        RECT 476.660 15.310 476.920 15.630 ;
        RECT 516.680 15.310 516.940 15.630 ;
        RECT 516.740 2.400 516.880 15.310 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 478.010 472.500 478.330 472.560 ;
        RECT 479.390 472.500 479.710 472.560 ;
        RECT 478.010 472.360 479.710 472.500 ;
        RECT 478.010 472.300 478.330 472.360 ;
        RECT 479.390 472.300 479.710 472.360 ;
        RECT 479.390 27.100 479.710 27.160 ;
        RECT 534.590 27.100 534.910 27.160 ;
        RECT 479.390 26.960 534.910 27.100 ;
        RECT 479.390 26.900 479.710 26.960 ;
        RECT 534.590 26.900 534.910 26.960 ;
      LAYER via ;
        RECT 478.040 472.300 478.300 472.560 ;
        RECT 479.420 472.300 479.680 472.560 ;
        RECT 479.420 26.900 479.680 27.160 ;
        RECT 534.620 26.900 534.880 27.160 ;
      LAYER met2 ;
        RECT 477.830 500.000 478.110 504.000 ;
        RECT 477.870 499.645 478.010 500.000 ;
        RECT 477.800 499.275 478.080 499.645 ;
        RECT 478.030 491.115 478.310 491.485 ;
        RECT 478.100 472.590 478.240 491.115 ;
        RECT 478.040 472.270 478.300 472.590 ;
        RECT 479.420 472.270 479.680 472.590 ;
        RECT 479.480 27.190 479.620 472.270 ;
        RECT 479.420 26.870 479.680 27.190 ;
        RECT 534.620 26.870 534.880 27.190 ;
        RECT 534.680 2.400 534.820 26.870 ;
        RECT 534.470 -4.800 535.030 2.400 ;
      LAYER via2 ;
        RECT 477.800 499.320 478.080 499.600 ;
        RECT 478.030 491.160 478.310 491.440 ;
      LAYER met3 ;
        RECT 477.775 499.620 478.105 499.625 ;
        RECT 477.750 499.610 478.130 499.620 ;
        RECT 477.750 499.310 478.560 499.610 ;
        RECT 477.750 499.300 478.130 499.310 ;
        RECT 477.775 499.295 478.105 499.300 ;
        RECT 478.005 491.460 478.335 491.465 ;
        RECT 477.750 491.450 478.335 491.460 ;
        RECT 477.750 491.150 478.560 491.450 ;
        RECT 477.750 491.140 478.335 491.150 ;
        RECT 478.005 491.135 478.335 491.140 ;
      LAYER via3 ;
        RECT 477.780 499.300 478.100 499.620 ;
        RECT 477.780 491.140 478.100 491.460 ;
      LAYER met4 ;
        RECT 477.775 499.295 478.105 499.625 ;
        RECT 477.790 491.465 478.090 499.295 ;
        RECT 477.775 491.135 478.105 491.465 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 480.310 26.420 480.630 26.480 ;
        RECT 552.530 26.420 552.850 26.480 ;
        RECT 480.310 26.280 552.850 26.420 ;
        RECT 480.310 26.220 480.630 26.280 ;
        RECT 552.530 26.220 552.850 26.280 ;
      LAYER via ;
        RECT 480.340 26.220 480.600 26.480 ;
        RECT 552.560 26.220 552.820 26.480 ;
      LAYER met2 ;
        RECT 479.210 500.000 479.490 504.000 ;
        RECT 479.250 499.360 479.390 500.000 ;
        RECT 479.250 499.220 479.620 499.360 ;
        RECT 479.480 483.070 479.620 499.220 ;
        RECT 479.480 482.930 480.540 483.070 ;
        RECT 480.400 26.510 480.540 482.930 ;
        RECT 480.340 26.190 480.600 26.510 ;
        RECT 552.560 26.190 552.820 26.510 ;
        RECT 552.620 2.400 552.760 26.190 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 480.540 499.160 480.860 499.420 ;
        RECT 480.630 498.340 480.770 499.160 ;
        RECT 481.230 498.340 481.550 498.400 ;
        RECT 480.630 498.200 481.550 498.340 ;
        RECT 481.230 498.140 481.550 498.200 ;
        RECT 481.230 483.720 481.550 483.780 ;
        RECT 481.230 483.580 495.260 483.720 ;
        RECT 481.230 483.520 481.550 483.580 ;
        RECT 495.120 483.440 495.260 483.580 ;
        RECT 495.030 483.180 495.350 483.440 ;
        RECT 495.030 20.640 495.350 20.700 ;
        RECT 570.010 20.640 570.330 20.700 ;
        RECT 495.030 20.500 570.330 20.640 ;
        RECT 495.030 20.440 495.350 20.500 ;
        RECT 570.010 20.440 570.330 20.500 ;
      LAYER via ;
        RECT 480.570 499.160 480.830 499.420 ;
        RECT 481.260 498.140 481.520 498.400 ;
        RECT 481.260 483.520 481.520 483.780 ;
        RECT 495.060 483.180 495.320 483.440 ;
        RECT 495.060 20.440 495.320 20.700 ;
        RECT 570.040 20.440 570.300 20.700 ;
      LAYER met2 ;
        RECT 480.590 500.000 480.870 504.000 ;
        RECT 480.630 499.450 480.770 500.000 ;
        RECT 480.570 499.130 480.830 499.450 ;
        RECT 481.260 498.110 481.520 498.430 ;
        RECT 481.320 483.810 481.460 498.110 ;
        RECT 481.260 483.490 481.520 483.810 ;
        RECT 495.060 483.150 495.320 483.470 ;
        RECT 495.120 20.730 495.260 483.150 ;
        RECT 495.060 20.410 495.320 20.730 ;
        RECT 570.040 20.410 570.300 20.730 ;
        RECT 570.100 2.400 570.240 20.410 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 498.250 17.580 498.570 17.640 ;
        RECT 587.950 17.580 588.270 17.640 ;
        RECT 498.250 17.440 588.270 17.580 ;
        RECT 498.250 17.380 498.570 17.440 ;
        RECT 587.950 17.380 588.270 17.440 ;
      LAYER via ;
        RECT 498.280 17.380 498.540 17.640 ;
        RECT 587.980 17.380 588.240 17.640 ;
      LAYER met2 ;
        RECT 481.970 500.000 482.250 504.000 ;
        RECT 482.010 498.340 482.150 500.000 ;
        RECT 482.010 498.200 482.380 498.340 ;
        RECT 482.240 484.005 482.380 498.200 ;
        RECT 482.170 483.635 482.450 484.005 ;
        RECT 498.270 25.995 498.550 26.365 ;
        RECT 498.340 17.670 498.480 25.995 ;
        RECT 498.280 17.350 498.540 17.670 ;
        RECT 587.980 17.350 588.240 17.670 ;
        RECT 588.040 2.400 588.180 17.350 ;
        RECT 587.830 -4.800 588.390 2.400 ;
      LAYER via2 ;
        RECT 482.170 483.680 482.450 483.960 ;
        RECT 498.270 26.040 498.550 26.320 ;
      LAYER met3 ;
        RECT 479.590 483.970 479.970 483.980 ;
        RECT 482.145 483.970 482.475 483.985 ;
        RECT 479.590 483.670 482.475 483.970 ;
        RECT 479.590 483.660 479.970 483.670 ;
        RECT 482.145 483.655 482.475 483.670 ;
        RECT 479.590 26.330 479.970 26.340 ;
        RECT 498.245 26.330 498.575 26.345 ;
        RECT 479.590 26.030 498.575 26.330 ;
        RECT 479.590 26.020 479.970 26.030 ;
        RECT 498.245 26.015 498.575 26.030 ;
      LAYER via3 ;
        RECT 479.620 483.660 479.940 483.980 ;
        RECT 479.620 26.020 479.940 26.340 ;
      LAYER met4 ;
        RECT 479.615 483.655 479.945 483.985 ;
        RECT 479.630 26.345 479.930 483.655 ;
        RECT 479.615 26.015 479.945 26.345 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 443.740 499.500 444.060 499.760 ;
        RECT 443.830 499.080 443.970 499.500 ;
        RECT 443.830 498.880 444.290 499.080 ;
        RECT 443.970 498.820 444.290 498.880 ;
        RECT 442.130 485.760 442.450 485.820 ;
        RECT 443.510 485.760 443.830 485.820 ;
        RECT 442.130 485.620 443.830 485.760 ;
        RECT 442.130 485.560 442.450 485.620 ;
        RECT 443.510 485.560 443.830 485.620 ;
        RECT 96.670 472.500 96.990 472.560 ;
        RECT 442.130 472.500 442.450 472.560 ;
        RECT 96.670 472.360 442.450 472.500 ;
        RECT 96.670 472.300 96.990 472.360 ;
        RECT 442.130 472.300 442.450 472.360 ;
      LAYER via ;
        RECT 443.770 499.500 444.030 499.760 ;
        RECT 444.000 498.820 444.260 499.080 ;
        RECT 442.160 485.560 442.420 485.820 ;
        RECT 443.540 485.560 443.800 485.820 ;
        RECT 96.700 472.300 96.960 472.560 ;
        RECT 442.160 472.300 442.420 472.560 ;
      LAYER met2 ;
        RECT 443.790 500.000 444.070 504.000 ;
        RECT 443.830 499.790 443.970 500.000 ;
        RECT 443.770 499.470 444.030 499.790 ;
        RECT 444.000 498.790 444.260 499.110 ;
        RECT 444.060 491.370 444.200 498.790 ;
        RECT 443.600 491.230 444.200 491.370 ;
        RECT 443.600 485.850 443.740 491.230 ;
        RECT 442.160 485.530 442.420 485.850 ;
        RECT 443.540 485.530 443.800 485.850 ;
        RECT 442.220 472.590 442.360 485.530 ;
        RECT 96.700 472.270 96.960 472.590 ;
        RECT 442.160 472.270 442.420 472.590 ;
        RECT 96.760 82.870 96.900 472.270 ;
        RECT 96.760 82.730 97.360 82.870 ;
        RECT 97.220 2.400 97.360 82.730 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 487.210 471.820 487.530 471.880 ;
        RECT 488.590 471.820 488.910 471.880 ;
        RECT 487.210 471.680 488.910 471.820 ;
        RECT 487.210 471.620 487.530 471.680 ;
        RECT 488.590 471.620 488.910 471.680 ;
        RECT 487.210 30.840 487.530 30.900 ;
        RECT 605.430 30.840 605.750 30.900 ;
        RECT 487.210 30.700 605.750 30.840 ;
        RECT 487.210 30.640 487.530 30.700 ;
        RECT 605.430 30.640 605.750 30.700 ;
      LAYER via ;
        RECT 487.240 471.620 487.500 471.880 ;
        RECT 488.620 471.620 488.880 471.880 ;
        RECT 487.240 30.640 487.500 30.900 ;
        RECT 605.460 30.640 605.720 30.900 ;
      LAYER met2 ;
        RECT 483.350 500.000 483.630 504.000 ;
        RECT 483.390 499.135 483.530 500.000 ;
        RECT 483.320 498.765 483.600 499.135 ;
        RECT 488.610 497.235 488.890 497.605 ;
        RECT 488.680 471.910 488.820 497.235 ;
        RECT 487.240 471.590 487.500 471.910 ;
        RECT 488.620 471.590 488.880 471.910 ;
        RECT 487.300 30.930 487.440 471.590 ;
        RECT 487.240 30.610 487.500 30.930 ;
        RECT 605.460 30.610 605.720 30.930 ;
        RECT 605.520 2.400 605.660 30.610 ;
        RECT 605.310 -4.800 605.870 2.400 ;
      LAYER via2 ;
        RECT 483.320 498.810 483.600 499.090 ;
        RECT 488.610 497.280 488.890 497.560 ;
      LAYER met3 ;
        RECT 483.295 498.785 483.625 499.115 ;
        RECT 483.310 497.570 483.610 498.785 ;
        RECT 488.585 497.570 488.915 497.585 ;
        RECT 483.310 497.270 488.915 497.570 ;
        RECT 488.585 497.255 488.915 497.270 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 514.810 17.240 515.130 17.300 ;
        RECT 623.370 17.240 623.690 17.300 ;
        RECT 514.810 17.100 623.690 17.240 ;
        RECT 514.810 17.040 515.130 17.100 ;
        RECT 623.370 17.040 623.690 17.100 ;
      LAYER via ;
        RECT 514.840 17.040 515.100 17.300 ;
        RECT 623.400 17.040 623.660 17.300 ;
      LAYER met2 ;
        RECT 484.730 500.000 485.010 504.000 ;
        RECT 484.770 499.815 484.910 500.000 ;
        RECT 484.700 499.445 484.980 499.815 ;
        RECT 516.210 488.395 516.490 488.765 ;
        RECT 516.280 448.570 516.420 488.395 ;
        RECT 515.360 448.430 516.420 448.570 ;
        RECT 515.360 420.970 515.500 448.430 ;
        RECT 514.900 420.830 515.500 420.970 ;
        RECT 514.900 17.330 515.040 420.830 ;
        RECT 514.840 17.010 515.100 17.330 ;
        RECT 623.400 17.010 623.660 17.330 ;
        RECT 623.460 2.400 623.600 17.010 ;
        RECT 623.250 -4.800 623.810 2.400 ;
      LAYER via2 ;
        RECT 484.700 499.490 484.980 499.770 ;
        RECT 516.210 488.440 516.490 488.720 ;
      LAYER met3 ;
        RECT 484.675 499.780 485.005 499.795 ;
        RECT 484.675 499.610 485.220 499.780 ;
        RECT 486.030 499.610 486.410 499.620 ;
        RECT 484.675 499.465 486.410 499.610 ;
        RECT 484.920 499.310 486.410 499.465 ;
        RECT 486.030 499.300 486.410 499.310 ;
        RECT 486.030 488.730 486.410 488.740 ;
        RECT 516.185 488.730 516.515 488.745 ;
        RECT 486.030 488.430 516.515 488.730 ;
        RECT 486.030 488.420 486.410 488.430 ;
        RECT 516.185 488.415 516.515 488.430 ;
      LAYER via3 ;
        RECT 486.060 499.300 486.380 499.620 ;
        RECT 486.060 488.420 486.380 488.740 ;
      LAYER met4 ;
        RECT 486.055 499.295 486.385 499.625 ;
        RECT 486.070 488.745 486.370 499.295 ;
        RECT 486.055 488.415 486.385 488.745 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 434.310 500.040 434.630 500.100 ;
        RECT 434.310 499.900 445.810 500.040 ;
        RECT 434.310 499.840 434.630 499.900 ;
        RECT 445.670 499.760 445.810 499.900 ;
        RECT 445.580 499.500 445.900 499.760 ;
        RECT 424.190 484.740 424.510 484.800 ;
        RECT 434.310 484.740 434.630 484.800 ;
        RECT 424.190 484.600 434.630 484.740 ;
        RECT 424.190 484.540 424.510 484.600 ;
        RECT 434.310 484.540 434.630 484.600 ;
        RECT 121.050 38.660 121.370 38.720 ;
        RECT 424.190 38.660 424.510 38.720 ;
        RECT 121.050 38.520 424.510 38.660 ;
        RECT 121.050 38.460 121.370 38.520 ;
        RECT 424.190 38.460 424.510 38.520 ;
      LAYER via ;
        RECT 434.340 499.840 434.600 500.100 ;
        RECT 445.610 499.500 445.870 499.760 ;
        RECT 424.220 484.540 424.480 484.800 ;
        RECT 434.340 484.540 434.600 484.800 ;
        RECT 121.080 38.460 121.340 38.720 ;
        RECT 424.220 38.460 424.480 38.720 ;
      LAYER met2 ;
        RECT 434.340 499.810 434.600 500.130 ;
        RECT 445.630 500.000 445.910 504.000 ;
        RECT 434.400 484.830 434.540 499.810 ;
        RECT 445.670 499.790 445.810 500.000 ;
        RECT 445.610 499.470 445.870 499.790 ;
        RECT 424.220 484.510 424.480 484.830 ;
        RECT 434.340 484.510 434.600 484.830 ;
        RECT 424.280 38.750 424.420 484.510 ;
        RECT 121.080 38.430 121.340 38.750 ;
        RECT 424.220 38.430 424.480 38.750 ;
        RECT 121.140 2.400 121.280 38.430 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 443.970 486.780 444.290 486.840 ;
        RECT 447.190 486.780 447.510 486.840 ;
        RECT 443.970 486.640 447.510 486.780 ;
        RECT 443.970 486.580 444.290 486.640 ;
        RECT 447.190 486.580 447.510 486.640 ;
        RECT 144.510 39.340 144.830 39.400 ;
        RECT 443.970 39.340 444.290 39.400 ;
        RECT 144.510 39.200 444.290 39.340 ;
        RECT 144.510 39.140 144.830 39.200 ;
        RECT 443.970 39.140 444.290 39.200 ;
      LAYER via ;
        RECT 444.000 486.580 444.260 486.840 ;
        RECT 447.220 486.580 447.480 486.840 ;
        RECT 144.540 39.140 144.800 39.400 ;
        RECT 444.000 39.140 444.260 39.400 ;
      LAYER met2 ;
        RECT 447.470 500.000 447.750 504.000 ;
        RECT 447.510 498.680 447.650 500.000 ;
        RECT 447.280 498.540 447.650 498.680 ;
        RECT 447.280 486.870 447.420 498.540 ;
        RECT 444.000 486.550 444.260 486.870 ;
        RECT 447.220 486.550 447.480 486.870 ;
        RECT 444.060 39.430 444.200 486.550 ;
        RECT 144.540 39.110 144.800 39.430 ;
        RECT 444.000 39.110 444.260 39.430 ;
        RECT 144.600 2.400 144.740 39.110 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 158.770 487.460 159.090 487.520 ;
        RECT 448.570 487.460 448.890 487.520 ;
        RECT 158.770 487.320 448.890 487.460 ;
        RECT 158.770 487.260 159.090 487.320 ;
        RECT 448.570 487.260 448.890 487.320 ;
      LAYER via ;
        RECT 158.800 487.260 159.060 487.520 ;
        RECT 448.600 487.260 448.860 487.520 ;
      LAYER met2 ;
        RECT 448.850 500.000 449.130 504.000 ;
        RECT 448.890 498.680 449.030 500.000 ;
        RECT 448.660 498.540 449.030 498.680 ;
        RECT 448.660 487.550 448.800 498.540 ;
        RECT 158.800 487.230 159.060 487.550 ;
        RECT 448.600 487.230 448.860 487.550 ;
        RECT 158.860 82.870 159.000 487.230 ;
        RECT 158.860 82.730 159.920 82.870 ;
        RECT 159.780 1.770 159.920 82.730 ;
        RECT 161.870 1.770 162.430 2.400 ;
        RECT 159.780 1.630 162.430 1.770 ;
        RECT 161.870 -4.800 162.430 1.630 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 450.180 499.500 450.500 499.760 ;
        RECT 445.350 497.660 445.670 497.720 ;
        RECT 450.270 497.660 450.410 499.500 ;
        RECT 445.350 497.520 450.410 497.660 ;
        RECT 445.350 497.460 445.670 497.520 ;
        RECT 179.930 39.680 180.250 39.740 ;
        RECT 445.350 39.680 445.670 39.740 ;
        RECT 179.930 39.540 445.670 39.680 ;
        RECT 179.930 39.480 180.250 39.540 ;
        RECT 445.350 39.480 445.670 39.540 ;
      LAYER via ;
        RECT 450.210 499.500 450.470 499.760 ;
        RECT 445.380 497.460 445.640 497.720 ;
        RECT 179.960 39.480 180.220 39.740 ;
        RECT 445.380 39.480 445.640 39.740 ;
      LAYER met2 ;
        RECT 450.230 500.000 450.510 504.000 ;
        RECT 450.270 499.790 450.410 500.000 ;
        RECT 450.210 499.470 450.470 499.790 ;
        RECT 445.380 497.430 445.640 497.750 ;
        RECT 445.440 39.770 445.580 497.430 ;
        RECT 179.960 39.450 180.220 39.770 ;
        RECT 445.380 39.450 445.640 39.770 ;
        RECT 180.020 2.400 180.160 39.450 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 451.560 498.820 451.880 499.080 ;
        RECT 451.650 498.340 451.790 498.820 ;
        RECT 451.650 498.200 452.020 498.340 ;
        RECT 450.870 497.660 451.190 497.720 ;
        RECT 451.880 497.660 452.020 498.200 ;
        RECT 450.870 497.520 452.020 497.660 ;
        RECT 450.870 497.460 451.190 497.520 ;
        RECT 450.870 488.480 451.190 488.540 ;
        RECT 427.730 488.340 451.190 488.480 ;
        RECT 193.270 488.140 193.590 488.200 ;
        RECT 427.730 488.140 427.870 488.340 ;
        RECT 450.870 488.280 451.190 488.340 ;
        RECT 193.270 488.000 427.870 488.140 ;
        RECT 193.270 487.940 193.590 488.000 ;
      LAYER via ;
        RECT 451.590 498.820 451.850 499.080 ;
        RECT 450.900 497.460 451.160 497.720 ;
        RECT 193.300 487.940 193.560 488.200 ;
        RECT 450.900 488.280 451.160 488.540 ;
      LAYER met2 ;
        RECT 451.610 500.000 451.890 504.000 ;
        RECT 451.650 499.110 451.790 500.000 ;
        RECT 451.590 498.790 451.850 499.110 ;
        RECT 450.900 497.430 451.160 497.750 ;
        RECT 450.960 488.570 451.100 497.430 ;
        RECT 450.900 488.250 451.160 488.570 ;
        RECT 193.300 487.910 193.560 488.230 ;
        RECT 193.360 82.870 193.500 487.910 ;
        RECT 193.360 82.730 195.800 82.870 ;
        RECT 195.660 1.770 195.800 82.730 ;
        RECT 197.750 1.770 198.310 2.400 ;
        RECT 195.660 1.630 198.310 1.770 ;
        RECT 197.750 -4.800 198.310 1.630 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 424.650 41.380 424.970 41.440 ;
        RECT 451.790 41.380 452.110 41.440 ;
        RECT 424.650 41.240 452.110 41.380 ;
        RECT 424.650 41.180 424.970 41.240 ;
        RECT 451.790 41.180 452.110 41.240 ;
        RECT 215.350 19.620 215.670 19.680 ;
        RECT 424.650 19.620 424.970 19.680 ;
        RECT 215.350 19.480 424.970 19.620 ;
        RECT 215.350 19.420 215.670 19.480 ;
        RECT 424.650 19.420 424.970 19.480 ;
      LAYER via ;
        RECT 424.680 41.180 424.940 41.440 ;
        RECT 451.820 41.180 452.080 41.440 ;
        RECT 215.380 19.420 215.640 19.680 ;
        RECT 424.680 19.420 424.940 19.680 ;
      LAYER met2 ;
        RECT 452.990 500.000 453.270 504.000 ;
        RECT 453.030 499.815 453.170 500.000 ;
        RECT 452.960 499.445 453.240 499.815 ;
        RECT 453.190 498.595 453.470 498.965 ;
        RECT 453.260 473.690 453.400 498.595 ;
        RECT 452.340 473.550 453.400 473.690 ;
        RECT 452.340 471.650 452.480 473.550 ;
        RECT 451.880 471.510 452.480 471.650 ;
        RECT 451.880 41.470 452.020 471.510 ;
        RECT 424.680 41.150 424.940 41.470 ;
        RECT 451.820 41.150 452.080 41.470 ;
        RECT 424.740 19.710 424.880 41.150 ;
        RECT 215.380 19.390 215.640 19.710 ;
        RECT 424.680 19.390 424.940 19.710 ;
        RECT 215.440 2.400 215.580 19.390 ;
        RECT 215.230 -4.800 215.790 2.400 ;
      LAYER via2 ;
        RECT 452.960 499.490 453.240 499.770 ;
        RECT 453.190 498.640 453.470 498.920 ;
      LAYER met3 ;
        RECT 452.935 499.465 453.265 499.795 ;
        RECT 452.950 498.945 453.250 499.465 ;
        RECT 452.950 498.630 453.495 498.945 ;
        RECT 453.165 498.615 453.495 498.630 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 454.320 499.700 454.640 499.760 ;
        RECT 454.320 499.500 454.780 499.700 ;
        RECT 439.830 496.980 440.150 497.040 ;
        RECT 454.640 496.980 454.780 499.500 ;
        RECT 439.830 496.840 454.780 496.980 ;
        RECT 439.830 496.780 440.150 496.840 ;
        RECT 227.770 488.820 228.090 488.880 ;
        RECT 439.830 488.820 440.150 488.880 ;
        RECT 227.770 488.680 440.150 488.820 ;
        RECT 227.770 488.620 228.090 488.680 ;
        RECT 439.830 488.620 440.150 488.680 ;
      LAYER via ;
        RECT 454.350 499.500 454.610 499.760 ;
        RECT 439.860 496.780 440.120 497.040 ;
        RECT 227.800 488.620 228.060 488.880 ;
        RECT 439.860 488.620 440.120 488.880 ;
      LAYER met2 ;
        RECT 454.370 500.000 454.650 504.000 ;
        RECT 454.410 499.790 454.550 500.000 ;
        RECT 454.350 499.470 454.610 499.790 ;
        RECT 439.860 496.750 440.120 497.070 ;
        RECT 439.920 488.910 440.060 496.750 ;
        RECT 227.800 488.590 228.060 488.910 ;
        RECT 439.860 488.590 440.120 488.910 ;
        RECT 227.860 82.870 228.000 488.590 ;
        RECT 227.860 82.730 233.520 82.870 ;
        RECT 233.380 2.400 233.520 82.730 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 440.520 499.360 440.840 499.420 ;
        RECT 440.520 499.220 441.440 499.360 ;
        RECT 440.520 499.160 440.840 499.220 ;
        RECT 441.300 498.060 441.440 499.220 ;
        RECT 441.210 497.800 441.530 498.060 ;
        RECT 55.730 479.640 56.050 479.700 ;
        RECT 441.210 479.640 441.530 479.700 ;
        RECT 55.730 479.500 441.530 479.640 ;
        RECT 55.730 479.440 56.050 479.500 ;
        RECT 441.210 479.440 441.530 479.500 ;
      LAYER via ;
        RECT 440.550 499.160 440.810 499.420 ;
        RECT 441.240 497.800 441.500 498.060 ;
        RECT 55.760 479.440 56.020 479.700 ;
        RECT 441.240 479.440 441.500 479.700 ;
      LAYER met2 ;
        RECT 440.570 500.000 440.850 504.000 ;
        RECT 440.610 499.450 440.750 500.000 ;
        RECT 440.550 499.130 440.810 499.450 ;
        RECT 441.240 497.770 441.500 498.090 ;
        RECT 441.300 479.730 441.440 497.770 ;
        RECT 55.760 479.410 56.020 479.730 ;
        RECT 441.240 479.410 441.500 479.730 ;
        RECT 55.820 2.400 55.960 479.410 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 75.970 486.780 76.290 486.840 ;
        RECT 442.130 486.780 442.450 486.840 ;
        RECT 75.970 486.640 442.450 486.780 ;
        RECT 75.970 486.580 76.290 486.640 ;
        RECT 442.130 486.580 442.450 486.640 ;
      LAYER via ;
        RECT 76.000 486.580 76.260 486.840 ;
        RECT 442.160 486.580 442.420 486.840 ;
      LAYER met2 ;
        RECT 442.410 500.000 442.690 504.000 ;
        RECT 442.450 498.680 442.590 500.000 ;
        RECT 442.220 498.540 442.590 498.680 ;
        RECT 442.220 486.870 442.360 498.540 ;
        RECT 76.000 486.550 76.260 486.870 ;
        RECT 442.160 486.550 442.420 486.870 ;
        RECT 76.060 82.870 76.200 486.550 ;
        RECT 76.060 82.730 79.880 82.870 ;
        RECT 79.740 2.400 79.880 82.730 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.110 18.940 103.430 19.000 ;
        RECT 445.810 18.940 446.130 19.000 ;
        RECT 103.110 18.800 446.130 18.940 ;
        RECT 103.110 18.740 103.430 18.800 ;
        RECT 445.810 18.740 446.130 18.800 ;
      LAYER via ;
        RECT 103.140 18.740 103.400 19.000 ;
        RECT 445.840 18.740 446.100 19.000 ;
      LAYER met2 ;
        RECT 444.250 500.000 444.530 504.000 ;
        RECT 444.290 499.815 444.430 500.000 ;
        RECT 444.220 499.445 444.500 499.815 ;
        RECT 445.830 498.595 446.110 498.965 ;
        RECT 445.900 19.030 446.040 498.595 ;
        RECT 103.140 18.710 103.400 19.030 ;
        RECT 445.840 18.710 446.100 19.030 ;
        RECT 103.200 2.400 103.340 18.710 ;
        RECT 102.990 -4.800 103.550 2.400 ;
      LAYER via2 ;
        RECT 444.220 499.490 444.500 499.770 ;
        RECT 445.830 498.640 446.110 498.920 ;
      LAYER met3 ;
        RECT 444.195 499.780 444.525 499.795 ;
        RECT 443.980 499.465 444.525 499.780 ;
        RECT 443.980 498.930 444.280 499.465 ;
        RECT 445.805 498.930 446.135 498.945 ;
        RECT 443.980 498.630 446.135 498.930 ;
        RECT 445.805 498.615 446.135 498.630 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 446.040 499.160 446.360 499.420 ;
        RECT 446.130 498.000 446.270 499.160 ;
        RECT 443.370 497.860 446.270 498.000 ;
        RECT 430.630 497.660 430.950 497.720 ;
        RECT 443.370 497.660 443.510 497.860 ;
        RECT 430.630 497.520 443.510 497.660 ;
        RECT 430.630 497.460 430.950 497.520 ;
        RECT 430.630 486.100 430.950 486.160 ;
        RECT 420.830 485.960 430.950 486.100 ;
        RECT 124.270 485.080 124.590 485.140 ;
        RECT 420.830 485.080 420.970 485.960 ;
        RECT 430.630 485.900 430.950 485.960 ;
        RECT 124.270 484.940 420.970 485.080 ;
        RECT 124.270 484.880 124.590 484.940 ;
      LAYER via ;
        RECT 446.070 499.160 446.330 499.420 ;
        RECT 430.660 497.460 430.920 497.720 ;
        RECT 124.300 484.880 124.560 485.140 ;
        RECT 430.660 485.900 430.920 486.160 ;
      LAYER met2 ;
        RECT 446.090 500.000 446.370 504.000 ;
        RECT 446.130 499.450 446.270 500.000 ;
        RECT 446.070 499.130 446.330 499.450 ;
        RECT 430.660 497.430 430.920 497.750 ;
        RECT 430.720 486.190 430.860 497.430 ;
        RECT 430.660 485.870 430.920 486.190 ;
        RECT 124.300 484.850 124.560 485.170 ;
        RECT 124.360 82.870 124.500 484.850 ;
        RECT 124.360 82.730 126.800 82.870 ;
        RECT 126.660 2.400 126.800 82.730 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 26.290 18.260 26.610 18.320 ;
        RECT 439.370 18.260 439.690 18.320 ;
        RECT 26.290 18.120 439.690 18.260 ;
        RECT 26.290 18.060 26.610 18.120 ;
        RECT 439.370 18.060 439.690 18.120 ;
      LAYER via ;
        RECT 26.320 18.060 26.580 18.320 ;
        RECT 439.400 18.060 439.660 18.320 ;
      LAYER met2 ;
        RECT 438.270 500.000 438.550 504.000 ;
        RECT 438.310 498.340 438.450 500.000 ;
        RECT 438.080 498.200 438.450 498.340 ;
        RECT 438.080 492.050 438.220 498.200 ;
        RECT 438.080 491.910 438.680 492.050 ;
        RECT 438.540 485.420 438.680 491.910 ;
        RECT 438.540 485.280 439.600 485.420 ;
        RECT 439.460 18.350 439.600 485.280 ;
        RECT 26.320 18.030 26.580 18.350 ;
        RECT 439.400 18.030 439.660 18.350 ;
        RECT 26.380 2.400 26.520 18.030 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.730 500.000 439.010 504.000 ;
        RECT 438.770 498.340 438.910 500.000 ;
        RECT 438.770 498.200 439.140 498.340 ;
        RECT 439.000 486.045 439.140 498.200 ;
        RECT 27.690 485.675 27.970 486.045 ;
        RECT 438.930 485.675 439.210 486.045 ;
        RECT 27.760 82.870 27.900 485.675 ;
        RECT 27.760 82.730 30.200 82.870 ;
        RECT 30.060 1.770 30.200 82.730 ;
        RECT 32.150 1.770 32.710 2.400 ;
        RECT 30.060 1.630 32.710 1.770 ;
        RECT 32.150 -4.800 32.710 1.630 ;
      LAYER via2 ;
        RECT 27.690 485.720 27.970 486.000 ;
        RECT 438.930 485.720 439.210 486.000 ;
      LAYER met3 ;
        RECT 27.665 486.010 27.995 486.025 ;
        RECT 438.905 486.010 439.235 486.025 ;
        RECT 27.665 485.710 439.235 486.010 ;
        RECT 27.665 485.695 27.995 485.710 ;
        RECT 438.905 485.695 439.235 485.710 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 405.330 784.185 694.590 787.015 ;
        RECT 405.330 778.745 694.590 781.575 ;
        RECT 405.330 773.305 694.590 776.135 ;
        RECT 405.330 767.865 694.590 770.695 ;
        RECT 405.330 762.425 694.590 765.255 ;
        RECT 405.330 756.985 694.590 759.815 ;
        RECT 405.330 751.545 694.590 754.375 ;
        RECT 405.330 746.105 694.590 748.935 ;
        RECT 405.330 740.665 694.590 743.495 ;
        RECT 405.330 735.225 694.590 738.055 ;
        RECT 405.330 729.785 694.590 732.615 ;
        RECT 405.330 724.345 694.590 727.175 ;
        RECT 405.330 718.905 694.590 721.735 ;
        RECT 405.330 713.465 694.590 716.295 ;
        RECT 405.330 708.025 694.590 710.855 ;
        RECT 405.330 702.585 694.590 705.415 ;
        RECT 405.330 697.145 694.590 699.975 ;
        RECT 405.330 691.705 694.590 694.535 ;
        RECT 405.330 686.265 694.590 689.095 ;
        RECT 405.330 680.825 694.590 683.655 ;
        RECT 405.330 675.385 694.590 678.215 ;
        RECT 405.330 669.945 694.590 672.775 ;
        RECT 405.330 664.505 694.590 667.335 ;
        RECT 405.330 659.065 694.590 661.895 ;
        RECT 405.330 653.625 694.590 656.455 ;
        RECT 405.330 648.185 694.590 651.015 ;
        RECT 405.330 642.745 694.590 645.575 ;
        RECT 405.330 637.305 694.590 640.135 ;
        RECT 405.330 631.865 694.590 634.695 ;
        RECT 405.330 626.425 694.590 629.255 ;
        RECT 405.330 620.985 694.590 623.815 ;
        RECT 405.330 615.545 694.590 618.375 ;
        RECT 405.330 610.105 694.590 612.935 ;
        RECT 405.330 604.665 694.590 607.495 ;
        RECT 405.330 599.225 694.590 602.055 ;
        RECT 405.330 593.785 694.590 596.615 ;
        RECT 405.330 588.345 694.590 591.175 ;
        RECT 405.330 582.905 694.590 585.735 ;
        RECT 405.330 577.465 694.590 580.295 ;
        RECT 405.330 572.025 694.590 574.855 ;
        RECT 405.330 566.585 694.590 569.415 ;
        RECT 405.330 561.145 694.590 563.975 ;
        RECT 405.330 555.705 694.590 558.535 ;
        RECT 405.330 550.265 694.590 553.095 ;
        RECT 405.330 544.825 694.590 547.655 ;
        RECT 405.330 539.385 694.590 542.215 ;
        RECT 405.330 533.945 694.590 536.775 ;
        RECT 405.330 528.505 694.590 531.335 ;
        RECT 405.330 523.065 694.590 525.895 ;
        RECT 405.330 517.625 694.590 520.455 ;
        RECT 405.330 512.185 694.590 515.015 ;
      LAYER li1 ;
        RECT 405.520 510.795 694.400 788.405 ;
      LAYER met1 ;
        RECT 405.520 510.640 694.400 788.560 ;
      LAYER met2 ;
        RECT 419.050 795.720 420.510 796.210 ;
        RECT 421.350 795.720 422.810 796.210 ;
        RECT 423.650 795.720 425.110 796.210 ;
        RECT 425.950 795.720 427.410 796.210 ;
        RECT 428.250 795.720 429.710 796.210 ;
        RECT 430.550 795.720 432.010 796.210 ;
        RECT 432.850 795.720 434.310 796.210 ;
        RECT 435.150 795.720 436.610 796.210 ;
        RECT 437.450 795.720 438.910 796.210 ;
        RECT 439.750 795.720 441.210 796.210 ;
        RECT 442.050 795.720 443.510 796.210 ;
        RECT 444.350 795.720 445.810 796.210 ;
        RECT 446.650 795.720 448.110 796.210 ;
        RECT 448.950 795.720 450.410 796.210 ;
        RECT 451.250 795.720 452.710 796.210 ;
        RECT 453.550 795.720 455.010 796.210 ;
        RECT 455.850 795.720 457.310 796.210 ;
        RECT 458.150 795.720 459.610 796.210 ;
        RECT 460.450 795.720 461.910 796.210 ;
        RECT 462.750 795.720 464.210 796.210 ;
        RECT 465.050 795.720 466.510 796.210 ;
        RECT 467.350 795.720 468.810 796.210 ;
        RECT 469.650 795.720 471.110 796.210 ;
        RECT 471.950 795.720 473.410 796.210 ;
        RECT 474.250 795.720 475.710 796.210 ;
        RECT 476.550 795.720 478.010 796.210 ;
        RECT 478.850 795.720 480.310 796.210 ;
        RECT 481.150 795.720 482.610 796.210 ;
        RECT 483.450 795.720 484.910 796.210 ;
        RECT 485.750 795.720 487.210 796.210 ;
        RECT 488.050 795.720 489.510 796.210 ;
        RECT 490.350 795.720 491.810 796.210 ;
        RECT 492.650 795.720 494.110 796.210 ;
        RECT 494.950 795.720 496.410 796.210 ;
        RECT 497.250 795.720 498.710 796.210 ;
        RECT 499.550 795.720 501.010 796.210 ;
        RECT 501.850 795.720 503.310 796.210 ;
        RECT 504.150 795.720 505.610 796.210 ;
        RECT 506.450 795.720 507.910 796.210 ;
        RECT 508.750 795.720 510.210 796.210 ;
        RECT 511.050 795.720 512.510 796.210 ;
        RECT 513.350 795.720 514.810 796.210 ;
        RECT 515.650 795.720 517.110 796.210 ;
        RECT 517.950 795.720 519.410 796.210 ;
        RECT 520.250 795.720 521.710 796.210 ;
        RECT 522.550 795.720 524.010 796.210 ;
        RECT 524.850 795.720 526.310 796.210 ;
        RECT 527.150 795.720 528.610 796.210 ;
        RECT 529.450 795.720 530.910 796.210 ;
        RECT 531.750 795.720 533.210 796.210 ;
        RECT 534.050 795.720 535.510 796.210 ;
        RECT 536.350 795.720 537.810 796.210 ;
        RECT 538.650 795.720 540.110 796.210 ;
        RECT 540.950 795.720 542.410 796.210 ;
        RECT 543.250 795.720 544.710 796.210 ;
        RECT 545.550 795.720 547.010 796.210 ;
        RECT 547.850 795.720 549.310 796.210 ;
        RECT 550.150 795.720 551.610 796.210 ;
        RECT 552.450 795.720 553.910 796.210 ;
        RECT 554.750 795.720 556.210 796.210 ;
        RECT 557.050 795.720 558.510 796.210 ;
        RECT 559.350 795.720 560.810 796.210 ;
        RECT 561.650 795.720 563.110 796.210 ;
        RECT 563.950 795.720 565.410 796.210 ;
        RECT 566.250 795.720 567.710 796.210 ;
        RECT 568.550 795.720 570.010 796.210 ;
        RECT 570.850 795.720 572.310 796.210 ;
        RECT 573.150 795.720 574.610 796.210 ;
        RECT 575.450 795.720 576.910 796.210 ;
        RECT 577.750 795.720 579.210 796.210 ;
        RECT 580.050 795.720 581.510 796.210 ;
        RECT 582.350 795.720 583.810 796.210 ;
        RECT 584.650 795.720 586.110 796.210 ;
        RECT 586.950 795.720 588.410 796.210 ;
        RECT 589.250 795.720 590.710 796.210 ;
        RECT 591.550 795.720 593.010 796.210 ;
        RECT 593.850 795.720 595.310 796.210 ;
        RECT 596.150 795.720 597.610 796.210 ;
        RECT 598.450 795.720 599.910 796.210 ;
        RECT 600.750 795.720 602.210 796.210 ;
        RECT 603.050 795.720 604.510 796.210 ;
        RECT 605.350 795.720 606.810 796.210 ;
        RECT 607.650 795.720 609.110 796.210 ;
        RECT 609.950 795.720 611.410 796.210 ;
        RECT 612.250 795.720 613.710 796.210 ;
        RECT 614.550 795.720 616.010 796.210 ;
        RECT 616.850 795.720 618.310 796.210 ;
        RECT 619.150 795.720 620.610 796.210 ;
        RECT 621.450 795.720 622.910 796.210 ;
        RECT 623.750 795.720 625.210 796.210 ;
        RECT 626.050 795.720 627.510 796.210 ;
        RECT 628.350 795.720 629.810 796.210 ;
        RECT 630.650 795.720 632.110 796.210 ;
        RECT 632.950 795.720 634.410 796.210 ;
        RECT 635.250 795.720 636.710 796.210 ;
        RECT 637.550 795.720 639.010 796.210 ;
        RECT 639.850 795.720 641.310 796.210 ;
        RECT 642.150 795.720 643.610 796.210 ;
        RECT 644.450 795.720 645.910 796.210 ;
        RECT 646.750 795.720 648.210 796.210 ;
        RECT 649.050 795.720 650.510 796.210 ;
        RECT 651.350 795.720 652.810 796.210 ;
        RECT 653.650 795.720 655.110 796.210 ;
        RECT 655.950 795.720 657.410 796.210 ;
        RECT 658.250 795.720 659.710 796.210 ;
        RECT 660.550 795.720 662.010 796.210 ;
        RECT 662.850 795.720 664.310 796.210 ;
        RECT 665.150 795.720 666.610 796.210 ;
        RECT 667.450 795.720 668.910 796.210 ;
        RECT 669.750 795.720 671.210 796.210 ;
        RECT 672.050 795.720 673.510 796.210 ;
        RECT 674.350 795.720 675.810 796.210 ;
        RECT 676.650 795.720 678.110 796.210 ;
        RECT 678.950 795.720 680.410 796.210 ;
        RECT 418.500 504.280 680.960 795.720 ;
        RECT 418.500 504.000 436.150 504.280 ;
        RECT 663.310 504.000 680.960 504.280 ;
      LAYER met3 ;
        RECT 421.050 510.715 663.055 788.485 ;
  END
END user_project_wrapper
END LIBRARY

